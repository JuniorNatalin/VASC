��   �*�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�NIO_AN_T�   L $�A* DR  �7SHIFT>V�ALID>I:I�E	IR�&CFG�.� �$V�ERSION �$COMME�NJ �USTOM� @ �2�DE_V_ENB> � �N�TMP�ST�ART_MODE~�NUM_LSJ��� �CHG_�DIG_PR�P�S_MAX���$� ;OP?] MKW>We�STr� ?I_OFS6O�] ��@q�����D<� KDV- KHO�L!�DH*ACT?_INDEX�c!�OPC�o!Kf*Kt)INIT�o �NNOT_NAM�� �$ORDE�= � �#HWl#�"R�EV�(SW1�*2r�*3#� SLO$�� VV3D 8IN��CP16XX_W&C51�D4��C53Y9PKX:PK~�SEARCH�� CHK�TP_�WA� c G�;M�AIN� Q>�2P�ARAM�7EXEyC6�R1SH2�S �HENABL�EpO^#SG_U}O�WD_TI� �;@ C� � P_DoEBUGPBSC,�?CS!DEFAUL�TPB�5�CAPD}U�PWRCLH<�1�KN_IO�A�K��!C�H�F�CFLA�G^#U!P�PWOFF_ALA� �BR� c"DBW@V��0�C.W�C�"2SY�;T[IO� �BOARD_S�!9B�T6�OP�YABD �XP�XMIS�U��W�ALM�Z�W��@`�U>A�Z� �YSM�VH�R� �XDc!iT�[�WmNOP fREAD�0�TS�T�D�fQ�1�j2�j3�UUP�DAT��0RC_�FIN@��aSI�Z�gJD�e>B�eDE��uPTH�fGR�OU��cOUJULONG�!Nt�!NtT1Nt4Kw5Kw6Kw�7Kw8KsBYTE �C�r�C�r1�tvq�t �q�t�q�t�q�t�q�tM9�w10��x1�x�1�x ��x1�x1��x1�x1�2����2. (d�f F)@�DI)0�ELTA#���	O�PT��W܆IOR_TRAN��ڄ�!RST�0��a��RESE�^PLI��1�S�"�INT#VL`L&X��O�!d�HO!$@ڀ�`@�ڀ�`@�U@RT�#���#��3�� vq���q���q���q�� �q���������(� ���@��ҙX���8p���FW_���1� 5 ��Wa�cN�CFIR�P@�W�\&DB. �{ �
BASE�V) � UsI��� vs��vs�료s���s�/�뢈���Y�T��6��~�y�Pb{���o � �RE�@p��>A!5LAYw���bt��}ADD �@�W��W�t3W� �T�5\�6\�7\�8���IA� �� ���!$CNaT��uP�6��RI����PROC�`���` ���`�źB�D ����0�#�5Ϙ|T�ǘ� A� �"X0���վ ��TYP������IP: < �����MAS�0��;pT�� ���QMSC�=�� �PrP>�Q�")�چ� O��"�D�!tF�UNK� �F��EXIl�C*`BUSY~���6*`�5��P� �槃@ B� U�Pr�F��FWV��SN��H���X1�`��� ��OCEX� A���� MAC��ML{FB��F_IP-����F_GW3�R3_1&U�U��SàCOU� �Ap�P1�� �� >AX3>A�>At3>Ay� >A��>A��>A��>A���� O�B��O���Z� ��e���p���{����s���s�USX3Oj� Pt3O��O��O��PO��O��(��L��� � $PA�TH_XDЀA ����	c�� 	c� (u#���N��E�� ����$DOWN�LOA�9@�ARAp܀�#M�" �����l u����ً������S�NU�K_��&�K8! B�OPER@�8�A��CHE��J!��D$	bhS%�#	cB:�	2A'CPYA%��#LO� ^&�11A'�1�O(SE�R&��A'P ���'��B!��&�&t1�(��eB�K$�@0BUP� Y�5R e&.6�2�'�#7�!7 �"���)���)���)����#�a_BT'#�2DTV�5���3�d�5�6 B!���C�5�C�5�s�5 �s�"�8��D��D�� ,D��@�'�RvG5P���BADb@�WNGsGS�G$�TIN:`N�EAFE��@_��&��LD�9I�A=���P���P��SERVLI,�(�h!o���{���#CM:WSVFZLOIW	b��fW��NR���'IO5��V곐�в�pU�U��"�~dMOn�b$H!CM� �S��b�@t�NY�e a#c�tet�.f+�D&d�CLzf0�_+���ID _� [�lge�lg o�lg��lg��lg��ްYNC_�vc�e�c �bsf�e�k�c�e�c�e��c�e�cHp� L�1v��C!C! �s!�s!�s!�s! �s!�s!�Nr�Nr|Rw(�CLASS��[����ve�����L�� 	 � >ΪENABL�����ES��+PENGTaHJ>��_�UB9������DA7�S�]��ϠR�ERRDEA�C�I#�NDEX ��3p���VPaQ�bh]��IM0x
� K$��H�"��L��ET���V��H�ٰ�bR5�0�BF��"I#�����R_Nv`P QIALB�$R7�0<Q1��_$VMA��MTSIMS��El��"� <���AƠ � 
Ϊ9���>�����PU%�摝�안� ��]�_�4����WRKxH 1v;v��	���`�0�"�\�TP_DEBUG�"гO�_�GPWO*0"�!W�  �a�Ns�������ɥ��OM����UBcYT�����$S_�SYSY����U�g�y��ϝ��$�s  ������Y�a �N��#AN 2 ���N� V�� ��Y����������ĵ˵Ա$�Ӳ��Ӳ�ӲI
-�ӲE�Ӳ]ϐӲ԰wϽ���Ӳ��Ӳ��Ӳ���Ͻ�I��Ӳ�ӲߒӲ 5�Ӳ"M�Ӳ$$e�Ӳ&}�Ӳ(��ӲI*��Ӳ,��Ӳ.���Ӳ0�߂��"CFG� ��V8�20P02 13O1028̵�����O�̵P��� :��� ~�Ӱ4�ś�@�����X��òX�FAN�UC Robot� Control�lerC�A05�B-2600-JS93 ��V|�� ?�  !�Y�V ��Y�d°������� ���ñ��U���, ���e�̵f�mc:�pniotrc.�txtX��ı��xX�������2 "�L�B�&А�N�C�y�İ�װ����)� �b�� 2��� hC�P1604 DA?P V2.6iђL�!"�X�#"�p�%$"���'"���5"��%7"�)"� �1°Lн� "�(M�̵������&�16�̲+= Oay��l��
�XX{ i���/"/�O/�/ �/�/�/?%?7?I? [???�?�?�?�?d����̲��?(O(O�?I��G ��;!� .1.��tM��1� �e���g�tO7OID����� �kjbv�tu211150�r01rs--kux�O	__-_?_Q_���V_z_�_�_�_�_��__WS7-PC �_oo,o>oPoboe_��o�o�o�o�o�o�j!�172.2d@8�.22hO�c255.&u�bw�V"�=Z~�c�� ����زj!'��l 6�Z�C�~�m�����Ə����ُ�V 	u�) ��!�Y��k�}�������ş�=L� ��AMC�:PCST_1.�X� ��+�AU�D1:\PN26�10.FWL 3�.9J�l+�i�̳�;Xd d�����������ʯܯ�  ��jo6�H�Z�l�~������7�FR:S7PRJ�ֿ�9����\fw_im?age.fwW�!��.�U�g�y��� G,X���s�|���@n ��ЂH��@��C����? x��e�e��r���EEE�G����(��z E(r��^!!�����7�d�r	y���ST' 2	�J��D{?5�?ސ�ߓ�p?���ׅ�������E��H �@;�!��K�5��Y�@s�!��*�����J���������L��a����	�!��"�D������s�v������£A�C���i������*����% � :��Wi��5�o��+=���|
��(3	��x���d �ZC�a�i�������E�/ ?A�x���%/C/	��Z(w/�/ ������8!/�/�/ ��(� �/T?f?F�x?�?�?}? �?�?�?�?O,O>OO bOtO�OUO�O�O�O�O �O_�O(_:_L__p_ �_�_c_�_�_�_�_ o o�_6oHoZo)o~o�o �oqo�o�o�o�o  �oDVh7��� �����.�� @�d�v�E��������� ���Տ*�<�N�� r���S�����̟��� ���8�J�\�+��� ��a���ȯگ����� "��F�X�j�9����� ����ֿ迷���0� ��T�f�x�GϜϮ��� ���������,�>�� b�t߆�Uߪ߼��ߝ� ������:�L��p� ���c������� � �$���H�Z�)�l��� ��q���������  2VhzI�� ����.@ dv�W��� ��/�*/</N// r/�/�/e/�/�/�/�/ ??�/8?J?\?+?�? �?�?s?�?�?�?�?O "O�?4OXOjO9O�O�O �O�O�O�O�O�O_0_ B__f_x_G_�_�_�_ �_�_�_o�_,o>oPo oto�oUo�o�o�o�o �o�o:L^- ���u��� � �$��H�Z�l�;��� ������؏ꏹ��� � 2��V�h�z�I����� �����
�ٟ.�@� �d�v���W�����Я �������<�N�� `�����e���̿޿�� ��&���J�\�n�=� �Ϥ�s������ϻ�� "�4��X�j�|�Kߠ� �߁����������0� B��f�x��Y���� ��������,�>�P� �t�����g������� ����(L^- ���u���� $6Zl;� ������� / 2/D//h/z/I/�/�/ �/�/�/�/
?�/.?@? R?!?v?�?�?i?�?�? �?�?OO�?<ONO`O /O�O�O�OwO�O�O�O �O_&_�OJ_\_n_=_ �_�_�_�_�_�_�_�_ "o4ooXojo|oKo�o �o�o�o�o�o�o0 BTx�Y�� ������>�P� b�1�����g���Ώ�� ����(���L�^�p� ?�����u���ܟ� �$�6��Z�l�~�M� ����Ư�����˯ � 2�D��h�z���[��� ¿Կ����
�ٿ�@� R�!�vψϚ�iϾ��� �ϱ���*���N�`� /߄ߖߨ�w������� ���&�8��\�n�=� ������������� "�4�F��j�|���]� ������������0 BT#x��k� ����>P b1���y�� ��/(/�L/^/p/ ?/�/�/�/�/�/�/ ? �/$?6??H?l?~?M? �?�?�?�?�?�?O�? 2ODOVO%OzO�O[O�O �O�O�O�O
__�O@_ R_d_3_�_�_i_�_�_ �_�_oo*o�_No`o roAo�o�o�o�o�o�o �o&8\n� O������� �4�F��j�|���]� ��ď֏������� B�T�#�x�����k��� ҟ䟳���,���P� b�1�t�����y�ί� ����(�:�	�^�p� ��Q�������ܿ� � Ͽ$�6�H��l�~ϐ� _ϴ��ϕ�������� 2�D�V�%�zߌߞ�m� �����ߵ�
����@� R�d�3����{��� �������*���<�`� r�A������������� ��&8Jn� O������ �4FX'|����$PNIO_I�M0 
�����N��k� V�A05B-�2600-J93�0eF174�606 ��k���LST 2�	�Dn;*�?�e�F'_$g|/K#�`R(�b/�/B+�$bY!�/�/�/��(Q�/�/
??Y%�Z/(8?�?L"�y4�j?|?�?"H!�4�#�!�?�O�;�!�1�/OO � J.H)?KO]O  �L.H�1�O�OA-�5�P�?�O%_L"�T�_(_i_"�[PBT�/[_m_ �6DEQ9O�_�_ ��X}O�_��_[�C�?po�_�UZolo~oj�o�o�o?��d�F_�oE�" �Q�1!q�?7I[s�Q !q�_{��]�� *��N�`�r�A����� ����ޏ���я&�8� �\�n���O�����ȟ ������ߟ4�F�� X�|���]���į֯�� �����B�T�f�5� ����k���ҿ俳�� �,���P�b�t�CϘ� ��yϼ��������(� :�	�^�p߂�Qߦ߸� �ߙ��� ���$�6�H� �l�~��_������ ������� �D�V�%� z�����m��������� 
.��Rd3� ��{���� *<`rA�� ����/�&/8/ J//n/�/�/a/�/�/ �/�/�/?�/4?F?X? '?|?�?�?o?�?�?�? �?OO�?BOTOfO5O �O�O�O}O�O�O�O�O _,_�OP_b_t_C_�_ �_�_�_�_�_o�_(o :o	oLopo�oQo�o�o �o�o�o �o6H Z)~�_��� ��� ��D�V�h� 7�����m���ԏ揵� 
��.���R�d�v�E� �����������ß� *�<��`�r���S��� ��̯����ѯ�8� J��n�����a���ȿ ڿ�����"��F�X� '�|ώϠ�o������� ����0���T�f�5� xߜ߮�}��������� �,�>��b�t��U� �����������(� :�L��p�����c��� ������ ��6H Z)~��q�� �� �DVh 7������ �/./�@/d/v/E/ �/�/�/�/�/�/?�/ *?<?N??r?�?S?�? �?�?�?�?OO�?8O JO\O+O�O�OaO�O�O �O�O�O_"_�OF_X_ j_9_�_�_�_�_�_�_ �_oo0o�_Tofoxo Go�o�o�o�o�o�o�o ,>bt�U �������� :�L��p�����c��� ʏ܏�� ��$��H� Z�)�l�����q�Ɵ؟ ꟹ�� �2��V�h� z�I������ԯ��� ǯ�.�@��d�v��� W�������п���տ *�<�N��rτϖ�e� �����ϭ�����8� J�\�+߀ߒߤ�s��� ���߻��"���4�X� j�9��������� �����0�B��f�x� G������������� ��,>Pt�U ������ :L^-���u ��� //$/�H/ Z/l/;/�/�/�/�/�/ �/�/�/ ?2??V?h? z?I?�?�?�?�?�?�? 
O�?.O@OOdOvO�O WO�O�O�O�O�O__ �O<_N__`_�_�_e_ �_�_�_�_oo&o�_ Jo\ono=o�o�oso�o �o�o�o"4X j|K����� ���0�B��f�x� ��Y�����ҏ����� ׏,�>�P��t����� g���Ο������� (�L�^�-�������u� ʯܯ��$�6�� Z�l�;���������ؿ ���˿ �2�D��h� z�Iόϰ��ϑ����� 
���.�@�R�!�v߈� ��i߾��ߟ����� ��<�N�`�/���� w���������&��� J�\�n�=��������� ��������"4X j|K����� ��0BTx �Y�����/ /�>/P/b/1/�/�/ g/�/�/�/�/??(? �/L?^?p???�?�?u? �?�?�?�?O$O6OO ZOlO~OMO�O�O�O�O �O�O�O _2_D__h_ z_�_[_�_�_�_�_�_�
on�$PNIO�_MOD 2����;aN��  @DAP V2.6o��Phdj`ka�_�SAFE 8 B�YTEzohc�hd{o32�o�V"hd7hc�fka �o~hdUa�d�b�as ^p�_����� ���$�6�	�Z�l� ?���������؏ꏽ� � �2��V�h�;�z� ������ԟ���˟��.��R�d�v�+gST�M  ;eNja+q����Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T��f�x���O_WR�K ;i ���_j�bC���}<��	�