��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �
  ����
��WVAMP_T �  $X�1  $X2�AY@��/FC~5  $2�ENBA $DTo  / _R2� d ENAB�LEDnSCHD�_NUMA ?��/ CFG5�� $GROUP��$z ACCEL�@�G$MAX�_FREQ�2 L��DWEL�DE�BUG�PREW�SOUT�P�ULSEASHsIFt 7TYP4�$USE_AE�F} 4$GDO��  f0 �r?�NpWE�AVE_TSK u�V�_GP��SUPPORT_�CFnCNVT_?DONE p }�k}GRP 2�r�� _� �}$� TIME1�to$2'EXT� �(1#&(MODE_�SW�CO3 SW�IT � `/ PH�AX6  4 �� ECC$�T�ERMNnPE�AKno!AL � \ � �!I֑$�!N_VSTAR�#!r"ؾ�"�%�CY�CL42 ��/ � Tv"b $�CUR_REL_܂ �! l/ WP�R5 � 
$wCEN� _RI3_RADIU��XIz ] ZI�MUTi!$ELEVATIONg5�� N�CONTI�NUOe2q �ME�XAC=PE�8��6  H~ ��UENCYA�I�TUD4�2RIG�HC�2LEBL_�ANG1 �O�TF_� 	��  $3A�bE�T��n3C!�$ORGjHFB)KjH��P��C�.�DLDW�HR�E�_�3�B�C��D�B�Cp�@�D�A�CCHG�G�	Q�F	Q�F	Q�FINC�G=Q�F=Q�F=Q�F؃AVCPYC� _T��\#�Y~P#�@SY��H)@�UPD�"0n�$$CL�ASS  �C���Q��8 �P�� �VA2�U��  ��?��@�  aa�U �To-o?oQoco�P�T�N 2 �[ �f��ue@O�i�oc�Q� � �U#a	`��`�d ��` �����=�������b ����.pqUcw- �ut(q��uvp�P�@�xu��d�aPq�h&�8���
�s,��!}a� u s�s�a�s��������֏b�Q�  �2�[
Ta�SI��}�v���F� ,�?1�' ��P�0��P�P�a�� 0�l�jk��ҟ������,�>�llFIGURE 8��3�:�a0�*�X�e� ۯү�������L��R�d�v������TOCIR1q�d ֿA���B�,�>���0�����:�`�B�����������nj� pq�(qG�V�E�@�����`+ݳ��� �ߩ߻���������x'�9�S�L��8%��B�5)��T� `���p���䏟�� w��#�5�G�Y�k�}����mkTrianglej���>� ,߂�L���D�Qc u������� �������X�+ X2D����� //'/9/�}, >l/�/���/? !?3?E?W?i?{?�?��C��?nhE��?�? OO,O>OPObOtO�O �O�O�O�O�O�K�?�O �?�?H_Z_l_~_�_�_ �_�_�_�_�_o o2o�|mSCHEXTENB  ��c��STATE 2�k @o�o�o�o��oNgWPR ����}��_OTOF 	�oa�@� �qq]qQcuv�quA��os�u@�  <#�
�?��^�1u�_GP 2;| �Io(�:���� ����e+