��   2W�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���C�ELL_GRP_�T   � �$'FRAME �$MOUN�T_LOCCCF�_METHOD � $CPY_SRC_IDX_�PLATFRM_�OFSCtDIM~_ $BASE{ �FSETC��A�UX_ORDER�   �X�YZ_MAP �� �LEN�GTH�TTCH�_GP_M~ a AUTORAIL_� �$$CLA�SS  ��i���D��D�8LOOR ���D8�?���O��/, � 1 F �H8=_`_��D'�82 �����K!/3/E//i/{/�-_ �/�/�/pO,��p 8!�/ �/?/g?y?�?]?�? �?�?�/�?�?�?�/C?E?�13OEOWOY?�O �O�O�O�O	__	O3_@E__1O�O�O�A{_ �_�_�O�_	oo�_?o�QocoQ_{o�ogo�$�MNU>A�R��d  8K=��q?�r�����?4ti���Ra?5}#?5�O�� ��4���D]  �P?��0��M �_=?Qs� �����	��� ?�)�K�u�_������� ���ˏ݋����ۏ 5�7�I�k������˟ ��ן���7�!�C� m�W�y�������ٯïկ����b!�K�2� G�i�k�}���ɿ��տ ����5��A�k�U� wϡϋϭ�������� ��	�C�-�?�a�c�u� ���߫��������-� �9�c�M�o���� ���������;�%�7�Y�[�A�1q����� ��������-9 cMo����� ��;%Gq [m������ �%//1/[/E/g/�/ {/�/�/�/�/�/�/	? 3????i?S?e?�?�?�?�?�?��A�?O�? O1O3OEOgO�O{O�O �O�O�O�O�O	_3__ ?_i_S_u_�_�_�_�_ �_�_o�_o)o+o=o _o�oso�o�o�o�o�o �o+7aKm ����������!�#�  �$M�NUFRAMEN_UM  W�>$��D  �k�TOOL A���������\ @�&�L����à?ϝ�D��Z�Ï3��S� 3��?�i�S�u����� ��՟�������A� +�=�_�a�s������� ˯��߯�+��7�a� K�m�������Ϳ��ٿ ����9�#�5�W�Y� kύϷϡ��������� #��/�Y�C�eߏ�y� ���߯���������1� �-�O�Q�c���� �����䲁p�����n� 2�4�F�h���|����� ��������
4@ jTv����� ���*,>` �t������ /,//8/b/L/n/�/ �/�/�/�/�/�/�/ ? "?$?6?X?�?l?�?�? �?�?�?�?�?$OO0O ZODOfO�OzO�O�O�O��O�O�O�O__
�1 3_q_X_m_�_�_�_�_ �_�_�_%oo1o[oEo go�o{o�o�o�o�o�o �o	3/iSe �������� �)�S�=�_���s��� ����ˏ��ߏ�+�� '�a�K�]�������� ߟɟ����!�K�5� W���k�������ï� ׯ��#���Y�C�U�w�y��A��Ϳ��ɿ ����!�K�5�Wρ� kύϷϡ��������� #��/�Y�C�eߏ�y� ���߯���������� C�-�O�y�c���� ����������'�Q� ;�]���q��������� ������;%Gq [}������ �I3Ui�{�����  ��$MNUTOO�LNUM  �
 
 D  @!