A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DMR_GRP_T  � $MASTER_DONE  $OT_MINUS   	$OT_PLUS   	$MASTER_COUN   	$REF_DONE  $REF_POS   	$REF_COUNT   	$BCKLSH_SIGN   	$EACHMST_DON   	$SPC_COUNT   	$SPC_MOVE   	$ADAPT_INER   	$ADAPT_FRIC   	$ADAPT_COL_P   	$ADAPT_COL_M   	$ADAPT_GRAV   	$SPC_ST_HIST   	$DSP_ST_HIST   	$SHIFT_ERROR  $SPC_CNT_HIS   	$MCH_PLS_HIS   	$ARM_PARAM   d$MASTER_ANG  $DSP_ST_HIS2   	$CLDET_CNT   	$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$GRAV_MAST   ��FMS_GRP_T t *$REM_LIFE   	$NT_LIFE   	$T_LIFE   	$CLDET_ANG   	$CLDET_DSTB   	$NT_LIFE_0   	$T_LIFE_TEMP   	$REM_LIFE_0   	$GRP_CL_TIME  $PCCOMER_CNT   	$FB_COMP_CNT   	$CMAL_DETECT   	$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $DTY_STR_T  $DTY_END_T  $CLDET_CNT   	$CLACT1   $CLACT2   $CLACT3   $CLACT4   $CLACT5   $CLACT6   $CL_OVR   $CLOMEGA1   $CLOMEGA2   $CLOMEGA3   $CLOMEGA4   $CLOMEGA5   $CLOMEGA6   $CL_FRMZ   $CLDEPT_IDX   $CLCURLINE   $CLDEST1   $CLDEST2   $CLDEST3   $CLDEST4   $CLDEST5   $CLDEST6   $CLNAME ?( �PLCL_GRP_T  � 	$CALIB_STAT  $TRQ_MGN   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	L�VCAX_REFA_T  @ $REF_FACTORY  $NUM_SET  $MAST_TO_REF  $PRE_MST2REF   ��VCAX_REFD_T  , $COMMENT $REF_UPDATE  $REF_AXIS 2 	H�VCAX_REFS_T  8 $STEP_MS_ENB  $NUM_SET  $STEP_DATA  $PRE_STEP  �VCAX_REFM_T   $IS_SET  $MASTER_COUN  �VCAX_REFG_T  0 $REF_DATA 2 
$REF_STEP 2 	$PRE_MASTER 2 	�$$CLASS  ������       �$DMR_GRP 1 ������      	                                      	                                      	 ��%��( �[�� [���                 	                                      	                                      	                                   	                                	 �dn� G �o{���xs6���             	                                      	                    	                    	                    	                    	 ���"�� J (       	                    	 B B B   B  B                   	 ���������K�_�����.��             	 ��#W��6����� [���             d                                                                                 =L��                                    ?�                              @�                                                                                                                                                                                                                                                           	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 �����$FMS_GRP 1������  	 I_t�H(�]IG�J<�J�>J.��             	 NdO¤*N�J:J�*sJ`��J(�             	 B�  B�  B�  B�  B�  B�               	 A�{CA�5��p�B�L��8���             	                                      	 Nt��P"�O0t�K�J�q�JN��             	 A�EA�EA�EA�EA�EA�E             	 I_v�H(��IG�|J<�J�uJ.�]            X�d 	                                      	                                      	                                                                V�|cV�vsV�V��WB/W��X�dN}��N}��N}�VN}�YN}�[Oi�COt�6Ou�R|u6S4XS4PV~wTV~ykX�Z�X�Z� 	    $                               ������8��ֱ���1������i��fF��rK d�y �� ��� ��.���f������}���b]��\~��V����7����  D�C�C�*C� C�eC��Z'E�' ��d�)�5�M�C��C�D)j�XC�~D�C�[Cߧ  ӕ��ȩѿ���ѡ�ѵ�N��"z��� �� ��� ����k�'�j�N��,[�4o����Ͳ  ��A����������D����/��I��`_T^5�����+��M�.����������  ���t��P��R���<���Z���Uj��T%����R ��`\(�`Z$�`W}��D���9���"7��n���5���3��H���I�  �����Fv��I���0,��SC��L���\���{��������������r��9���,������cD��(��$���>���>�        d   d   d   d   d   (   
   (   (   (   (   d   d   d   d   d   d   d   d  ����                                        ��������            s      ����    ����    ��������       ����       ����           ����������������  ����       ����    ����                             ����                ����      ����   ����                                       ����                         ����            ����                   ����        ����������������          ����                    ������������            ����   ��������   ����     e   e   e   e   e   e   e   e   e   e   e   e   e   e   e   e   e   e   e   e                            9                                                         "                  (      8   A   A   A            $   S   S   /   /  >Q�>P|>O��>P��>O�e>O�>�`8>T󘾵�f��oپ�P���X>PR�>P�N>QX >�`8>PŲ>Pڜ>P3d>PC�  ?Z�R?ZJ�?ZFR?Zj.?Z8�?ZA�?X?[~ž!M�>�&�>�4�>�X�?Z\�?Zn�?Z��?X?Zum?Zy�?ZU�?ZW�  �wkr�z���z���zH��z���z����w��{���@K����� ���zi��z=ھy�Ⱦ�w��z-x�z"��zz�z�?  <��<��w<���<��<���<���?�81<�+�?8���%���&���)<��v<���<��?�81<��]<��<��*<��{  ���Ϳ�ڿ�p��$���>���������?��f�$��$�_�$�c�� y��&��2�����(8��)���]��K  ?���?��B?���?���?���?��y�	��?����p��59�59��59�?���?��[?��)�	��?��o?���?���?���  ,($UP021                                     ($UP001...........................0050      ($UP001...........................0050      ($UP001...........................0050      ($UP001...........................0050      ($UP001...........................0050      ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001...........................0050      ($UP001...........................0050      ($UP001...........................0050      ($UP001                                     ($MAKRO080                                  ($MAKRO080                                  ($MAKRO080                                  ($MAKRO080                                   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      �$PLCL_GRP 1������� D    	 ?�  ?�  ?�  ?�  ?a]?s{?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$VCAX_REF_GR 2������ t 
 �REFERENCE 1        	                                                                                                                                                 REFERENCE 2        	                                                                                                                                                 REFERENCE 3        	                                                                                                                                                 REFERENCE 4        	                                                                                                                                                 REFERENCE 5        	                                                                                                                                                 REFERENCE 6        	                                                                                                                                                 REFERENCE 7        	                                                                                                                                                 REFERENCE 8        	                                                                                                                                                 REFERENCE 9        	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE2_1       	                                                                                                                                                 REFERENCE2_2       	                                                                                                                                                 REFERENCE2_3       	                                                                                                                                                 REFERENCE2_4       	                                                                                                                                                 REFERENCE2_5       	                                                                                                                                                 REFERENCE2_6       	                                                                                                                                                 REFERENCE2_7       	                                                                                                                                                 REFERENCE2_8       	                                                                                                                                                 REFERENCE2_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE3_1       	                                                                                                                                                 REFERENCE3_2       	                                                                                                                                                 REFERENCE3_3       	                                                                                                                                                 REFERENCE3_4       	                                                                                                                                                 REFERENCE3_5       	                                                                                                                                                 REFERENCE3_6       	                                                                                                                                                 REFERENCE3_7       	                                                                                                                                                 REFERENCE3_8       	                                                                                                                                                 REFERENCE3_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE4_1       	                                                                                                                                                 REFERENCE4_2       	                                                                                                                                                 REFERENCE4_3       	                                                                                                                                                 REFERENCE4_4       	                                                                                                                                                 REFERENCE4_5       	                                                                                                                                                 REFERENCE4_6       	                                                                                                                                                 REFERENCE4_7       	                                                                                                                                                 REFERENCE4_8       	                                                                                                                                                 REFERENCE4_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                         