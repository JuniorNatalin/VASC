��    ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�NSF_SET_�T   h �$MODE  �$IN_SIZ�<OUTDADD�RESS=BY_�PWFAIL= �fLCCONpR�U}T1ONLY�p`�$$CLA~`  ����:��U��U�$'1 ��U���������