��   t��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���U�I_CONFIG�_T  d �9$NUM_MENUS  9�* NECTCRE�COVER>CCOLOR_CRR�:EXTSTAT���$TOP>_�IDXCMEM_�LIMIR$D�BGLVL�PO�PUP_MASK��zA  $DUMMY54��ODE�
5CFO�CA �6CPS�)C��g HA�N� � TIME�OU�PIPES�IZE � MW�IN�PANEM;AP�  � � �FAVB ?� 
w$HL�_DIQ�?� qELEM�Z�UR� l� S|s�$HMI��RO+\W AD�ONLY� �T�OUCH�PRO�OMMO#?$��ALAR< �F�ILVEW�	E�NB=%%fC �1"USER:)FC[TN:)WI�� I* _ED�l"V!�_TITL� ~1"COORDF<#/LOCK6%�$F%|�!b"EBFOR�? �"e&
�"�%�!�BA�!j ?�"B�G�%$PM�X�_PKT�"IHE�LP� MER�B�LNK$=ENAB��!? SIPMAN�UA�-4"="�B�EEY?$�=&q!E�Dy#x&UST�OM0 t �$} RT_SPI�D��4C�4*PA�G� ?^DEV�ICE�9SCREVuEF���7N��@$FLAG�@�,�&�1  h� 	$PWD_A�CCES� E �8��TC�!�%)$�LABE� 	$	Tz j4@q!�D��	?\&USRV�I 1  < �`� �B��APRI�m� U1�@�TRIP�"m�$�$CLA?@ �����A��R��R��$'2 ~����R�	 �,��?���/Q�>P8R3T.Q��|��)P� UPyU_��
 ���A��_�_�_�_�_�_o  �_*o<oNo`oro�oo �o�o�o�o�o�o&�8J\n���(�/SOFTP�0/�GENLINK?�current=�menupage?,935,1�� ���!:�L�^�p� ����#���ʏ܏� � ���6�H�Z�l�~��� ��1�Ɵ؟���� � ��D�V�h�z�������� TPT�X����:�ٯ�� �s Ƿ���$/�softpart�/genlink�?help=/m�d/tp�q.dg@��F�X�j�|�5�&�#�pwd2�ɿۿ� ��4�#�5�G�Y�k�}� ϡϳ��������ϊ� ��1�C�U�g�yߋ�aT���AsVQR�� ($ ����������(����A2QN�PS�2S�������^�
�q�2QVQ��RQ  ���ʡ��	���E�����L�L�Y�9S�2 1�E>P�R \ }|mPREG �VED��6�H�w�holemod.�htm\�sing}lm�doub���trip��?brows���� I�������3EW�i{�3�W�i�d/ev.sr�l���	1�	t ��	 ��o��]��p���(/� �@ @/R/d/v/�/�/�/�/�/�/�& @</?#? �/G?Y?k?:6+�#// �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O��O�O#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo go5/�o�o�o�o�o�o  2D??hzI [��y?�?qo
�� �)�R�M�_�q����� �����ݏ��*�%� 7�_W�Q�������� ǟٟ����!�3�E� W�i�{�������ï�o ���"�4�F�X�j�|� �����Ŀֿ����� ���ͯf�a�sυ� �ϩϻ��������� >�9�K�]߆߁ߓ�a� �߭��������#�5� G�Y�k�}������ ���������Z�l� ~��������������� �� 2hz1� C�)�����
 )RM_q�� �������/	/ 7/I/[/m//�/�/�/ �/�/�/�/?!?3?E? W?i?{?I��?�?�?�? �?O"O4OFOXOS|O��O]OoO�O�O�J�$�UI_TOPME?NU 1�@Q�R 
�XQ�1)*de�fault�?�=	�*level0; *HP 8_& �o__m_Rtpi�o[23](tpst[1�X�_�_��_BVX_�_!$
h5�8e01.gif�o(	menu5Bi9`da13BjcbAjbad4ikPoa���o �o�o $6�2�o�_q����Ht�prim=dapa�ge,1422,1����/�A�L�e�w���������N���vclass,5�ȏ���!�3�E�P�܌13L���������4ʟQ��|53����*�<�N�Q��|8 ����������ѯP���@��+�=�O��9P Q_��B]y�aw��o�ÿ�Vty�]�_�Qm�f[0�_��	�c�[164�W>�59@�Xa�oٿ{�]h2�o gm��}j�osgAk���c g�y�F�X�j�|ߎ�� ������������0�B�T�f�x���ۍ2 ������������� O�a�s�����&�8�p�������� ۟�1�4�^p���%�~�sainedi����%�wintp�p0bt� ���6Qr���f o��//0/B/T/f/ x/�/ o�/�/�/�/�/ ??,?>?c?�o�?�? �?�?�?�? �OO)O ;OMO_O�?�O�O�O�O �O�O�O~O_%_7_I_ [_m_�O�_�_�_�_�_ �_z_o!o3oEoWoio {o
o�o�o�o�o�o�o �o/ASew ��������o�0������⯿]?o��s󽌏������u��d�f���&�4�Ӡ��B�h��ό�6��u7���0����'� 9��]�o��������� F�ۯ����#�5�G�
64�1C������� ��ɿԯ����#�5� G�ֿk�}Ϗϡϳ��� ��2�����1�C�U�����6\ߑߣߵ�����4Ӝ74��'� 9�K�]�������/ z����������"�G� F���R�|��������� ������p?1CUg y�Vϯ���� 	�?Qcu� �(����// �;/M/_/q/�/�/�/ 6/�/�/�/??%?�/ I?[?m??�?�?2?�? �?�?�?O!O3O�?WO iO{O�O�O�Ol�~��O ��l�
_._@_R_w_ v_�_�__�_�_�_o oo*o<oNo�o�o �o�o�o�o�oHO' 9K]o�o��� ���|�#�5�G� Y�k�}������ŏ׏ ������1�C�U�g� y��������ӟ��� 	���-�?�Q�c�u��� �����ϯ����O �O;��O�_^op����� ����ʿܿ�\���7� 6�H�Z�l�~ϐϢ�po �������!�3�Eߜ� i�{ߍߟ߱���R��� ����/�A�S���w� �������`���� �+�=�O���s����� ��������n�' 9K]������ ��j�#5G Yk&����ϲ�� ���//0/B/� b/`/�/�/�/�/�/�/ �/?��??Q?c?u?�? �?��?�?�?�?OO �?;OMO_OqO�O�O�O 6O�O�O�O__%_�O I_[_m__�_�_2_�_ �_�_�_o!o3o�_Wo io{o�o�o�o@o�o�o �o/�oSew ����z��� ??*�<�N�`�r��� �������ޏ���� &�K�J�\�*?������ ɟ۟�D�#�5�G� Y�k�}������ůׯ ������1�C�U�g� y��������ӿ��� 	Ϙ�-�?�Q�c�uχ� ϫϽ�������ߔ� )�;�M�_�q߃ߕ�$� �����������w�t�*defaul�t�w�*level8ˏi�{��7�� tpst[�1]����y��t?pio[23�����u��n��6�H�	�menu7.gi5fI�
h�13m�z��5��g��e�4��u6m�����%7 I��m���� V��!3EW~�prim=h��page,74,1\�������pclass,13�/(/:/L/^/��5d/�/�/�/�/�/���/?.?@?0R?d?gy18��?@�?�?�?�?�/�6�?�%O7OIO[OmOL��$�UI_USERV?IEW 1�q�q�R 
��tON�O�OF�m�O__%_7_I_�O m__�_�_�_X_�_�_ �_o!o�O.o@oRo�_ �o�o�o�o�oxo�o /AS�ow�� ��jo���b+� =�O�a�s�������� ͏ߏ����'�9�K�~�*zoom^�ZOOM]���� ԟ���
���.�@� R�d�v��������Я����*max�res��MAXRES������\�n� ������G�ȿڿ��� ϳ�4�F�X�j�|�'� �ϛϭ�������� 0�B���f�xߊߜ߮� Q�����������'� =�K�߆������ q�����(�:�L��� p���������c����� ��[�$6HZl �����{�  2D��Ucu� �����
/�./ @/R/d/v//�/�/�/ �/�/��/??�/N? `?r?�?�?9?�?�?�? �?OO�?8OJO\OnO �O#A