A��*SYSTEM*   V8.2306       4/24/2014 A5  *SYSTEM*  ��AAVM_WRK_T  � $EXPOSURE  $CAMCLBDATE $PS_TRGVT   $TRGVT  $TRGHZ  $TRGDIST  $TRGW  $TRGP  $TRGR  $LENS_CENT_X  $LENS_CENT_Y  $DISTORT   $CMP_GC_P  $UTNUM  $PRE_MAST_CT   	$PRE_GRV_MST  $NEW_MAST_CT   	$NEW_GRV_MST  $STAT_RUN  $RES_ERR  $VTCP_ERR   $TRGT_ERR   $RES_ERR2  $VTCP_ERR2   $RSM_MAST_CT   	$STAT_START  $STAT_END  $STAT_ORGBK  $STAT_RSMBK  $STAT_ORGRES  $STAT_UPDT  �ABSPOS_GRP_T   $PARAM    ��ALRM_RECOV_T    $ALMRECOVENB   $ALMRECOVON   �ALMDG_T  0 $DEBUG1  $DEBUG2  $DEBUG3  $CONT_TYPE  �ALM_IF_T  D $ENABLE  $LAST_ALM d$LAST_UALM d$KALM_MAX  $LDEBUG   
  ��APCOUPLED_T  $ $APP_PROCES0  $APP_PROCES1    D�APCUREQ_T  � $SOFTPART_ID  $TOTAL_EQ  $CUR_EQNO  $PS_SPI_INDE   $SPI_INDEX  $SCREEN_NAME $APP_SIGN $APP_PROCES0  $APP_PROCES1  $TOPK_FILE 	$THKY_FILE 	$PANE_EQNO   	$DUMMY12  $DUMMY13  $DUMMY14  @�ARG_STR_T  � $TITLE $ITEM1 $ITEM2 $ITEM3 $ITEM4 $ITEM5 $ITEM6 $ITEM7 $ITEM8 $ITEM9 $ITEM10 $ITEM11 $ITEM12 $ITEM13 $ITEM14 $ITEM15 $ITEM16 $ITEM17 $ITEM18 $ITEM19 $ITEM20 8�ASBN_CFG_T  8 $CNV_JNT_POS  $DATA_CMNTS  $FLAGS   $POS_CHECK  �AT_CELLSETUP 	 P $HOME_IO_PRG %$HOME_MACRO %$REPR_MACRO %$PRODRUN_SPD  $PRODRSM_SPD  D�AUTOBACKUP_T 
 $ENABLE  $DEVICE $TIME   $DI_IDX  $STARTUP_BCK  $INTERVAL  $DISP_UNIT  $BCK_DO_IDX  $ERR_DO_IDX  $FR_FREE  $IN_PROGRESS  $REQ_BACKUP  $PRC_WAIT  $AUTO_BACKUP  $POFF_COUNT  $DEL_COUNT  $LOG_IDX  $DEL_TIME ? $DEL_FILE ?� $PROC_FILE �@�MOTOR_COUNTE  0 $REM_COUNTS   	$REM_REV   	$BIL_REV   	 �AXIS_COUNTER   $ODOMETER $NON_CMD  D�AXIS_METER_T    $ODOMETER   	$NON_CMD   	 ��AXSCRDCFG_T  d $CARD_EXIST  $FSSB_TYPE  $CHKBD_SEL  $DIAG_REG   $SLOT_NUM  $SLOT_PREV  $DEBUG    ��BACK_EDIT_T  � $PROGRAM %$SRC_NAME %$EPT_IDX  $OPEN_ID  $DELETE_OK  $USED_TP_CRT  $BACKUP_NAME %$PS_REPLACIN   $REPLACING  $BCK_COMMENT $D_REPLACING  $SEL_PROGRAM %$DUMMY12  $DUMMY13  8�BLAL_OUT_T  , $DO_INDEX  $PS_BATALM_O   $BATALM_OR  �CFCFG_T  X $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $COMP_SWITCH  $MAX_NSETS  �CF_PARAMGP_T  � 
$WARNMESSENB  $CHKJNTLIM  $CNSTNT_CORN  $TIMEFLTRENB  $TRATIO_TB   $ACCTIME_TB1   $ACCTIME_TB2   $ORIENT_TYPE  $DEBUG  $RTSPD_SF   ��CHG_PRI_T   $TASK_ID  $PRIORITY   @�CHKPOS_T  x $CONT_FLAG  $POS_HDR  $JPOS1  $JPOS2  $JPOS3  $JPOS4  $JPOS5  $JPOS6  $JPOS7  $JPOS8  $JPOS9    ��COCFG_T  < $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $ENABLED  �CO_MORGRP_T  t $FLEN  $ANGLE  $TBA_MAG  $TBA_MAG_PRE  $TBA_MAG_MAX  $TBA_MAGAXS   	$TBA_CURAXS   	$TBA_PRVAXS   	H�CO_PARAMGP_T  � $OPT_TIME  $OPT_ACC  $JACC_RRATIO  $CACC_RRATIO  $JTIME_RATIO  $CTIME_RATIO  $JVARDMAX  $CVARDMAX  $WARNMESSENB  $DEBUG  $TBA_MGN  @�CP_RSMOFST_T  @ $RO_ENABLE  $RO_MAX_ITP  $RO_NOM_DIST  $RO_NOM_SPD   �CPCFG_T  � $GROUP_MASK  $CP_DEBUG  $CP_ENABLE  $COMP_SWITCH  $EXTRA_INT   $EXTRA_FLT   
$TF_MODE  $MD3ITPTOL  $RESUME_OFST $CP_HSTART  $T1_HSTART  $TEST   $COMP_SW2  $COMP_SW3  $COMP_SW4  �CPDBGDEF_T  d $OUTPUT  $FILENAME )$GROUP_MASK  $DEBUGMASK  $MAXDATA  $COUNT  $TAIL  $BUFEXIST  �CPDBG_T  � $OUTPUT  $CPIDEBUG $CPPDEBUG $MIDEBUG $MPDEBUG $MGDEBUG $MFDEBUG $SIMQSTOP  $KEEP  $PATH )$EXTRA1  $EXTRA2  �CP_L64FIX_T  � $ENABLE  $DEC_A   $DEC_V   $DEC_CIF   $DEC_PCHO   $ADD_A   $ADD_V   $ADD_CIF   $ADD_PCHO   $DEBUG_SIM  $SIM_ADDRESS  $SIM_VAR_TYP  $SIM_AXIS  $EXTRA1  $EXTRA2  $EXTRA3  �CP_MCRGRP_T  4 $RSM_JBF_PCT  $RSM_DEC_PCT  $RSM_OFS_PCT   ,�CP_MORGRP_T  � $CHNS_EMPTY  $GTF_EMPTY  $CHK_T1_SPD  $T1_FPSPD  $T1_TCPSPD  $SPEED  $T1SPDLIM  $SPEEDTOL  $JNT_VEL   	$JNT_ACC   	$JNT_JRK   	$SEGFRACTION  $RSTRT_LINE  $RSTRT_PVF  D�CP_TESTDEF_T    $ENABLE_TEST  $NUM_LINES  D�CP_PARAMGP_T  D )$WARNMESSENB  $DEBUG  $ENB  $NUM_CHN  $NUM_JBFSET  $NUM_JBF  $EXT_NUM_JBF  $JBF_SIZE  $EXT_JBF_SIZ  $NUM_TF  $TF_SIZE  $EXT_TF_SIZE  $NUM_RSINFO  $JNT_VEL_LIM   	$JNT_ACC_LIM   	$JNT_JRK_LIM   	$T1SEGFL_SF  $T1GTFL_SF  $CRCMP_SWITC  $ACCLIM_SF  $JRKLIM_SF  $PSPD_SWITCH  $MAX_PSPD  $MIN_PSPD  $PSPDACC_SF  $PSPDJRK_SF  $CDCOMP_SW  $CDACC_SF  $CDJRK_SF  $CDDELTATOL  $CDDISTSF  $CDANGTOL  $CDDEVTOL  $CHKJNTLIM  $FDANG_TOL  $FDLIN_TOL  $JNTJBF_ENB  $COMP_SW  $EXTRA_INT   $EXTRA_FLT   $CP_TEST H�CP_T1_MODE_T ! � 	$ENABLE  $COMP_SWITCH  $MARGIN  $TIME_FACTOR  $SPD_LIMIT  $SLEW_RATE  $MIN_TFLEN  $EXTRA_INT   $EXTRA_FLT     ��CRCFG_T "� $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $PGDEBUG  $CR_ENHANCED  $LGORN_ENBL  $BLEND_ENB  $MAX_ARC_ANG  $RSM_RSPD_LM  $LGORN_METH  $LGORN_DBG  $LGORN_RAD  $LGORN_AZ_SP  $LGORN_ELTOL  $ROTSPDFCTR  $MAX_FP_SPD  $SMCRC_RADI  $SMCRC_RADO  $SMCRC_ARC  $ARCANGLIM  $MAXORNTCHG  $MAXSGRATIO  $CHKBMP  $RSM_TYP  $CHK_MSK  $AES_SINGTOL  ��CRI_CFG_T #  $CRI_SW  �CSXC_PARAM_T $ x 	$NAME $ATTR  $NUM_CHANNEL  $IMG_HEIGHT  $IMG_WIDTH  $VT_SPACING  $DEF_ASPECT  $MIN_EXPO  $MAX_EXPO  �CUSTOMMENU_T % $ $TITLE $PROG_NAME %$OPTION  �CZ_CDCFG_T & x $ENABLE   $CD_ENABLE  $NO_HEADER  $COMP_SWITCH  $WARNMESSENB  $EXTRA_INT   $EXTRA_FLT   $CHK_SPD_SF  ��DBPXWORK_T '  $SKP_DEL   �DBTB_CTRL_T ( � $ACRT_MODE  $MINDT_ADJ  $DELAY_CALL  $DELAY_DO  $DELAY_PLS  $RESERVED1  $RESERVED2  $RESERVED3  $NUM_IO  $DUMMY9  $DUMMY10  d�DB_DBG_T )  $DBG_PRM   
��DPOS_DAT_T *  $X  $Y  $Z  �LDPOS_DAT_T +  $X  $Y  $Z  ��PD_T ,  $X  $Y  $Z  �PC_T -  $X  $Y  $Z  P�PENETRATE_T .  $X  $Y  $Z   �DB_RECORD_T /H $CPOS *$LPOS +$DPOS_DST  $LDPOS_DST  $LINE_NUM  $ONCE_DC  $CROSS  $TASK_ID  $ENABLED_TIM  $TRIGGER_TIM  $PAUSED_TIME  $RETURNED_TI  $MMR_STATUS $CRE_NEWMON  $SIGNAL_ACT  $LAST_ACT  $PD ,$PC -$PN_AT .$PD2  $PC2  $PT  $PD_DOT_PC  $LINE_DST  $P_NUM  $GO_AWAY  $MOTION_COMP  �DCSS_DEVICE_ 0 P $TYPE  $RBT_NUM  $SPI_IDX  $SPO_IDX  $SPI_BYTE  $SPO_BYTE  $STO  �DCSS_LS_T 1 H $STOOUT_IDX  $STOFB_IDX  $STOFB_CH  $FENCE_TYPE  $FENCE_IDX  �DCSS_PARAM_T 2 H $DOCHK_ENB  $PMCS_ENB  $LS_STOP  $LS_FENCE  $HOTSWP_TIME    ��DCSS_ELEM_T 3 T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    �DCSS_RBT_T 4 � $MDL_ELEM 23 
$ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$FB_TOL   	$RBT_TYPE  �DCS_CFG_T 5� $DISP_MENU  $LOG_ENB  $LOG_LEN  $LOG_FILE $LOG_ID  $LOG_IDMAX  $LOG_DELAY  $LOG_WRT  $LOG_INTVL  $LOG_EVENT  $TEST_PARAM1  $TEST_PARAM2  $CHK_J_TOL  $CHK_C_TOL  $SAFE_SPD  $SAFE_SPD_SV  $EXCLUDE   $SPD_ONLY   $SYS_PARAM  $PROTECT  $HI_VRC  $APPLY_WARN  $HIDE_MENU  $HI_VRC_MLT   $VRFY_ALL  $HI_MATE  $IOC_PROT  $IOC_CRC1  $IOC_CRC2  $OPI_VRC  �DCS_CRC_OUT_ 6  $START_GRP    �DCS_SGN_T 7 � 
$CURR_SIGNAT  $CURR_DATE $PREV_SIGNAT  $PREV_DATE $ANNUNC_TYP  $ANNUNC_IDX  $CUR_TIME   $LATCH_TIME   $CUR_CRC   $LATCH_CRC    �DEFLOGIC_T 8 @ $FUNC_TITLE 	$TOTAL_NUM  $DUMMY2  $DUMMY3  $DUMMY4  �DEMO_INIT_T 9 L $DEMO_ENB  $DEMO_AU  $DEMO_DAYS  $LOAD_NUM  $DUMMY4  $DUMMY5  �EFF_AXIS_T :  $NUM  $COEFF  �ADJ_RTRQ_T ; D $COR_TRQ   $COR_TEMP   $EFF_AXIS 2: $LIMIT  $ADJ_NUM  �AMP_COEF_T < 0 $COEF_A   	$COEF_C  $MASK  $DUAL_MASK  �CTRL_CAB_T = @ $TRANS_A  $IDLE_PWR  $AMP_COEFB  $SV_NUM  $SV_AMP 2< �DIAG_GRP_T >8 *$VAL_SET  $TACC   	$TACC_LIM1   	$TACC_LIM2   	$RRATE_LOAD   	$VER $ANSWER  $RCC_ANS  $ADJ_RTRQ 2; $ADJ_OHTRQ   	$COPPER   	$IRON   	$BRK_PWR   	$CABLE_ACT   $CABLE_BASE   	$CABLE_LENG   	$CAB_NUM  $CTRL_CAB 2= $TRQCNS   	$TRQDWN   	$MSBAS   	$MAXTRQ   	$RRATE   	$LIFECALC   	$L10   	$N0   	$T0   	$CUR_L10   	$TCP_TYPE  $CUR_TCP $MOTN_STYLE  $FLAG  $CUR_OVC   	$CUR_HEAT   	$SUPPORT_TYP   	$ALL_SUPPORT  $CUR_TCP_X  $CUR_TCP_Y  $CUR_TCP_Z  $CUR_TCP_W  $CUR_TCP_P  $CUR_TCP_R  �h�DICT_CFG_T ? ` $CACHE_ENB  $CACHE_SIZE  $CURR_ONLY  $LANG_SUFFIX $LOCALE  $DUMMY5  $DUMMY6   	��DMSW_CFG_T @ 8 $KEYIMAGE  $TMS_DSB  $TMS_STAT  $TMS_INPUT    �DOCVIEWER_T A  $DBGLVL  $CURFILE ?� 	p�DPM_CFG_T B x 
$ENABLE  $DPM_INLINE  $GRP_MSK  $BEF_JBF  $DELAY  $ORI_CTL  $CUR_SCH  $MAX_SCH  $COMP_SW  $DEBUG  ��OFS_CHN_T C � $ENABLE  $OTF_DI_IDX  $CHN_TYP  $RAMP_GAIN  $SCAN_RATE  $INI_OFS  $REM_OFS  $APP_OFS  $IN_TICK  $OU_TICK  $ID  $STAT  $MAX_LIM  $MIN_LIM  $MAX_INC  $MIN_INC  $A1  $A2   ��AI_CHN_T D  $P_GAIN  $D_GAIN  $I_GAIN  $STR_CNT  $REF_CNT  $AVE_CNT  $FBK_MODE  $REF_VAL  $RAW_FBK  $CAL_FBK  $PORT_NUM  $CAL_DONE  $SLOPE  $INTERCEPT  $CUR_TICK  $LEAD_DIS  $BUF_SIZE  $BUF_CNT  $T_ADJ  $MIN_VAL  $MAX_VAL  7��BI_CHN_T E D $DI_IDX1  $DI_IDX2  $BUMP_OFS  $BUMP_RATE  $BUMP_GAIN  t�GI_CHN_T F  $DI_IDX  $SCALE  (�DPM_GRP_T G � $OFS_TYPE  $OFS_FRAM  $LAST_DPM  $OFS_ACCU  $OFS_ABS  $OFS_CARRY  $CTL_RATE  $INT_LINE  $OFS_LINE  $DAT_RDY  $OFS_STAT  $SND_TYPE  $TRK_MODE  $SYNC_DI  $OFS 2C 	$AI_CH 2D 	$BI_CH 2E 	$GI_CH 2F 	��DPM_SCH_T H 0 $GRP_MSK  $COMMENT $DPM_ON  $GRP 2G '��DPM_IN_T I 8 $LINE_NUM  $DELAY  $OFS_X  $OFS_Y  $OFS_Z  ��DRC_CFG_T J D $HOST1 !$HOST2 !$HOST3 !$HOST4 !$HOST5 !$EMAIL_ENABL  ��DSBL_FAULT_T K  $ENABLE  $MAX_COUNT  ��DTREC_T L, $DTREC_ENB  $SAMPLE_ITP  $BUF_SIZE  $FILE_SIZE  $DEVICE_NAM $SUBBUF_SIZ  $SPC_FILE  $DTREC_ON  $DTSAV_ON  $FILE_ACCESS  $PC_ACCESS  $SYSTIME   P$DTSAV_ENB  $ORDER  $DSB_BUFSIZ  $ENB_BUFSIZ  $OTTASK_MOD  $DP_ALM_ID  $DP_ALM_GRP  $DP_ALM_AXS  $DEF_MAXBUF  ��DYN_BRK_T M 0 $DI_IDX  $DO_IDX  $BRK_MSK  $FLTR_IF  ��ENC_STAT_T N� $ENC_COUNT  $ENC_ROS_TIK  $ENC_RATE  $ENC_AVERAGE  $ENC_ENABLE  $ENC_DSPSTAT  $ENC_SPCSTAT  $ENC_SIM_ON  $ENC_SIM_SPD  $ENC_VALUE  $ENC_HEAD  $ENC_MULTIPL  $ENC_STOPPED   $ENC_THRESH  $ENC_EXISTS  $ENC_HSDI  $ENC_ABSCNT  $INCTRAVDIST  $INCTRAVCNTS  $INCTRAV_DO  $CONVSPD_GO  $INCTRAVRES  $ENC_BUFFER   d$ENC_ATR_AXS  $SC_GRP_NUM  $ENC_COMERCT  $ENC_FBCMPCT  �ENETMODE_T O 8 $FULL_DUPLEX  $SPEED  $ACD_ENABLE  $THROTTLE  <�ER_NOAUTO_T P D $NOAUTO_ENB  $NOAUTO_NUM  $PS_NOAUTO_C   $NOAUTO_CODE    H�ER_NOALM_T QH *$NOALMENBLE  $NOALM_NUM  $ER_CODE1  $ER_CODE2  $ER_CODE3  $ER_CODE4  $ER_CODE5  $ER_CODE6  $ER_CODE7  $ER_CODE8  $ER_CODE9  $ER_CODE10  $ER_CODE11  $ER_CODE12  $ER_CODE13  $ER_CODE14  $ER_CODE15  $ER_CODE16  $ER_CODE17  $ER_CODE18  $ER_CODE19  $ER_CODE20  $ER_CODE21  $ER_CODE22  $ER_CODE23  $ER_CODE24  $ER_CODE25  $ER_CODE26  $ER_CODE27  $ER_CODE28  $ER_CODE29  $ER_CODE30  $ER_CODE31  $ER_CODE32  $ER_CODE33  $ER_CODE34  $ER_CODE35  $ER_CODE36  $ER_CODE37  $ER_CODE38  $ER_CODE39  $ER_CODE40  Z��ER_OUTPUT_T R � $OUT_NUM  $IN_NUM  $PLCWARN  $GRP_STR  $ERROR_NUM  $FAC_NUM  $SEV_NUM  $PARM1_NUM  $PARM2_NUM  $DUMMY9  $DUMMY10  $DUMMY11   ��EXT_SET_T S < $ENABLE  $DI_TYPE  $DI_NUM  $DO_TYPE  $DO_NUM  �FDR_GRP_T TT $VEL_MOD   	$VEL_CNT   	$REM_LIFE2   	$OVM_RATE   	$OVA_RATE   	$TROV_RATE   	$DTAV_RATE   	$DTMX_RATE   	$DTMIN_RATE   	$MOT_RATE   	$DIAG_INDX_R   
$DIAG_INDX_I   $DG_MAXT   	$DG_T0   	$RATED_TRQ   	$DRIVE_TYPE   	$GEAR_RATIO2   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$Z_MCMD   	��FEATURE_T U , $NAM ? $MOD ? $VER ? $MEC ?  p�FILECOMP_T V  $TPP  $VARIABLE  ��FILE_SETUP2_ W 4 $FILE_TDC_SC  $FILE_TV_SEC  $FILE_TVC_SC   �FILE_BACK_T X T $FILE_NAME )$PROG_NAME %$FUNC_CODE  $MODIFIER  $COMMENT %$FUNC_PTR   ��FMR2_GRP_T Y $VEL_ROT  $VEL_LIN  $VEL_MOD   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$TROV_MAX   	$T_LIFE_0  $RATED_TRQ   	$LIMIT_FUNC  $ACC_LMT   	$DRIVE_TYPE   	$GEAR_RATIO2   	$DGCLFR   	$DGDYFR   	$DGLDEC   	$DG5T0   	$DG_MAXT   	$DG_T0   	��FMR_CFG_T Z  $TROV_MAX   T�FSSB_CFG_T [ P $FSSB_LINE   $EX_FSSBLINE   $FSSB1_AXES  $FSSB3_AXES  $FSSB5_AXES  �GRAVC_GRP_T \ � 
$MODE_SW  $SPCONS   	$DEBUG1  $DEBUG2   	$GRV_STATUS  $BKUP_NO116   	$POFF_NO116   	$GRVCMP_SW  $GRVMST_LOOP  $MST_SMT_LEN   H�MOTYPE_E ]       �TERMTYPE_E ^      �ORIENT_E _    a M�SM_PROFILE_E `    X���TA_PROFILE_E a       �UPR_T b� -$MOTYPE ]$TERMTYPE ^$SEGTERMTYPE ^$DECELTOL  $USE_CONFIG  $USE_TURNS  $ORIENT_TYPE _$UFRAME $UTOOL $SPEED  $ROTSPEED  $CONTAXISVEL  $CNSTNT_PATH  $CNSTNTPTHJT  $SEG_TIME  $USE_CARTACC  $USEMAXACCEL  $USERELACCEL  $USETIMESHFT   $USE_PATHACC  $USE_SHORTMO  $SM_PROFILE  `$TA_PROFILE  a$ACCEL_OVRD  $TIME_SHIFT  $ACCU_NUM   $PAYLOAD  $DYN_I_COMP  $PATHRES_ENB  $RESERVE1   $CNT_SHORTMO  $EXT_SPEED  $CNT_ACCEL1  $CNT_ACCEL2  $CRCCOMPENB  $ASYMFLTRENB  $USE_WJTURNS  $EXT_INDEP  $CARTFLTRENB  $CNT_SPEEDUP  $CNT_DYN_ACC  $MAX_SPEED  $USERELPSPD  $PSPD_OVRD  $ORNT_MROT  H�GRSMT_GRP_T c  $GRV_SW  $GRV_PARAM  d�HOST_CFG_T d � $COMMENT $PROTOCOL 	$PORT $OPER  $STATE  $MODE $REMOTE $REPERRS  $TIMEOUT  $PATH e$STRT_PATH e$STRT_REMOTE $USERNAME e$PWRD_TIMOUT  $SERVER_PORT  $USE_VIS_PRT  ��HOSTENT_T e 4 $H_NAME !$H_ADDRTYPE  $H_LENGTH  $H_ADDR !��ERR_MASK_T f H $SSC_MASK1  $SSC_MASK2  $SSC_MASK3  $SSC_MASK4  $SEV_MASK  4�HSCD_MNG_T g $COLL_MODE  $THRESHOLD  $DO_ERR  $DO_ENABLE  $MACRO_REG  $STND_CD  $AUTO_RESET  $UPD_GROUPS  $PARAM_VERID 	$PARAM119   	$PARAM120   	$PARAM121   	$PARAM122   	$PARAM123   	$PARAM124   	$PARAM125   	$ACT_RATIO  $SAVED119   	$SAVED120   	��HSCD_GRP_T h $ $COL_DET_OFF  $HSCD_PRM_ID   �HTTP_AUTH_T i ( $OBJECT !$NAME $TYPE  $LEVEL  �HTTP_T j � $ENABLE  $ENAB_DIAGTP  $ENAB_SPART  $DBGLVL  $KRL_TIMOUT  $HITCOUNT  $BG_COLOR $ENAB_TEMPL  $TEMPLATE $COMMENT $RSS_INUM  �HWR_CONFIG_T k H $MAINCPU  $VISIONCPU  $SPARE1  $SPARE2  $SPARE3  $SPARE4  ��IBGN_CFG_T l $CMP_WAIT  $MAX_PNUM1  $MAX_PNUM2  $FWD_TOL_LOC  $FWD_TOL_ORT  $FWD_TOL_EXT  $FWD_TOL_ANG  $BWD_TOL_LOC  $BWD_TOL_ORT  $BWD_TOL_EXT  $BWD_TOL_ANG  $BWD_RTN_SPD  $UF_DATA  $DBG_MASK  $TEMP_MGN  $LIN_N_CNST  $END_TOL_LOC  $STATUS  $RECDAT_SEND  ��IBGN_ERRIO_T m @ $REC_IO_TYP  $REC_IO_NUM  $EXE_IO_TYP  $EXE_IO_NUM   ��IBGN_EXEC_T n ( $SCHEDULE   $FILE_P   $BWD_FLG    ��IBGN_FIL_T o @ $EXE_MD  $EXE_OPN  $EXE_BACK  $REC_TRANS  $REC_ACC  �IBGN_FTP_T px $FTP_CTAG  $AUTO_TRANS  $IGNR_COMER  $FTP_STAG  $SM_STAG  $SM_CTAG  $SM_SPORT  $SM_CPORT  $N_PCSOFT 	$N_RECFL1 	$N_RECFL2 	$N_RECFL3 	$N_EXEFIL $N_FLEXT1 $N_CONDFL 	$N_FLEXT2 $N_SPTXT1 $N_SPTXT2 	$SEQ_VAR  $SNS_NUM  $SNS_CNST  $FOLDER $RECS_PRG %$RECS_TMO  $RECE_PRG %$RECE_TMO  $SM_DBG  $AUTO_START  $RESERVE  ��IOLNK_T q 8 $RACK  $SLOT  $INPUT_N  $OUTPUT_N  $OPTION   �IOSLAVE_T r  $INPUT_N  $OUTPUT_N  8�IO_DEF_ASG_T s T $LOG_TYPE  $LOG_NO  $NUM_PORTS  $RACK  $SLOT  $PHY_TYPE  $PHY_NO   �IO_UOP_CFG_T t ` $UOP_TYPE  $IN_RACK  $IN_SLOT  $IN_STRTPT  $OUT_RACK  $OUT_SLOT  $OUT_STRTPT   8�UJR_GRP_T u � $FINE_OVRD  $JOGFRAME $FINE_DIST  $J7_GROUP  $J8_GROUP  $J7_AXIS  $J8_AXIS  $J7_LABEL $J8_LABEL $J7_GRAPHIC Q$J8_GRAPHIC Q$DSB_J7J8  $DSBL_KEY   �KAREL_CFG_T v 0 $CONV_ENABLE  $CONV_CTRL  $CONV_FLAGS   ��LGCFG_T w � $ENABLE  $OUT_SW  $LG_SIZE  $EV_SIZE  $MR_SIZE  $SG_SIZE  $FD_SIZE  $MI_SIZE  $ER_SIZE  $MP_SIZE  $MG_SIZE  $PE_SIZE  $LG_MODE  $EV_MODE  $MR_MODE  $SG_MODE  $FD_MODE  $PE_MODE  $EX_RSCH_FIL $COMP_SW  ��LN_DISP_T x ` $HIDE_LINE_N  $DISP_MENU  $HIDE_PARLN  $HIDE_DAULN  $HEAD_PARENT $HEAD_DAUGHT  ��LOGBOOK_T yt B$NUM_ER_ITM  $NUM_ER_TYP  $NUM_REC_TYP  $NUM_SCRN_FL  $NUM_DIO  $SRAM_MARGIN  $DRAM_MARGIN  $OPTION  $LOG_ER  $LOG_ENT  $LOG_SEL  $LOG_WIN  $LOG_MENU  $LOG_JGMU  $LOG_MNCHG  $LOG_FNKEY  $LOG_JGKY  $LOG_PRGKEY  $LOG_UFKY  $LOG_OVRKY  $LOG_FWDKY  $LOG_HLDKY  $LOG_STPKY  $LOG_PRVKY  $LOG_ENTKY  $LOG_ITMKY  $LOG_RSTKY  $LOG_HELPKY  $LOG_OVR  $LOG_CRD  $LOG_STEP  $LOG_GRP  $LOG_SGRP  $LOG_UF  $LOG_UT  $LOG_FILE  $LOG_WTRLS  $LOG_PGCHG  $LOG_SETPOS  $LOG_TPKY  $LOG_DIO  $LOG_STMD  $LOG_FOCUS  $LOG_PRGEXE  $LOG_TUIKEY  $IMG_ENT  $IMG_SEL  $IMG_WIN  $IMG_FNKY  $SAVE_FILE 	$SCRN_FL  $SCRN_NO_ENT  $ANALOG_TOL  $AVAILABLE  $CLEAR_ENB  $DCS_HI1  $DCS_HI2  $DCS_HO1  $DCS_HO2  $DCS_SI  $DCS_SO1  $DCS_SO2  $DCS_OPTION  $IGNR_SAVE  $FNKEY_FLTR  $DCS_DEV  H�LOG_BUFF_T z 0 $TITLE $SIZE  $MEM_TYPE  $VISIBLE   ��LOG_STAT_T { 0 $TICK  $SPD  $POS1  $POS2  $POS3   ��LOG_DCS_T | � $ENABLE  $SPD_TOL  $OUTPUT_TYP  $OUTPUT_IDX  $GRP_NUM  $POS_TYP  $AXIS_NUM  $STOP_READY  $STOP {$ESTOP {$CSTOP {$ESTOP_DIFF {$CSTOP_DIFF { `�LOG_DIO_T } L $RACK  $SLOT  $MOD_TYPE  $PORT_TYPE  $START_PORT  $END_PORT   ��LOG_SCRN_FL_ ~  $SP_ID  $SCRN_ID  p�MCSP_T  � $CLDPOP_ENB  $TRQLIM_ENB  $JOGLIM_ENB  $CLDPOP_FLG  $CLDGRP_FLG  $CLDREL_FLG  $CLR_CLDFLG  $JOGLIM_FLG  $ORGJOG_OVR  $COMP_SW  $RESERVE1  $RESERVE2  $RESERVE3  \�MCSP_GRP_T � � 	$JOGLIM_OVR  $TRQLIM_FLG  $SV_PTLIM   	$ORG_PTLIM   	$ORG_RCLMC   	$RESERVE1  $RESERVE2  $RESERVE3   	$RESERVE4   	��MISC_GRP_T � d $HPD_TRQ   	$DSTB_MAX   	$DSTB_MIN   	$DSTB_MAXENB   	$DSTB_MINENB   	$DSTB_EXCESS   T�MISC_MSTR_T �  $HPD_ENB   h�MISC_SCD_T � H $DSTB_MAX_A   	$DSTB_MIN_A   	$DSTB_MAXENB   	$DSTB_MINENB   	��MKCFG_T � \ $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $MO_CONFLICT  $MO_REQUIRED  $DEBUG  l�MLTARM_CFG_T �  $NUM_ARMS  $GROUP   d�MLT_GRP_DO_T � � $TP_ENABLE  $JOG_GROUP  $LOCKED_ARM  $CRNT_TYPE  $CRNT_INDX  $PRG_ROUT_P  $JOG_ROUT_P  $PRG_DO_TYPE   $PRG_DO_INDX   $JOG_DO_TYPE   $JOG_DO_INDX    ��MNDSP_MST_T � ` $DISP_ENABLE  $DISP_EDCMD  $DISP_INAUTO  $DISP_RSMDIS  $DISP_IS_ON  $MODE_GRP   ��MNDSPPSTL_T � 4 $LOCTOL  $ORIENTTOL  $EXTTOL  $ANGTOL   	l�MODAQ_CFG_T � d $ON_LINE  $MF_FLAG  $MI_FLAG  $GRP_NUM  $STARTLOG  $ENDLOG  $LN_MASK  $SUPPORT   ��FX_TRIGGER_T � � 	$START_MODEL  $START_STEP  $START_PROG %$STOP_MODEL  $STOP_STEP  $STOP_PROG %$AXES  $DATA_TYPE  $DATETIME  �MODEM_INF_T � t $MDM_INIT )$MDM_INIT1 )$MDM_RESET )$MDM_HANGUP )$MDM_DIAL )$MDM_ANSWER )$MDM_STATUS )$MDM_IDENT )��MOR_GRP_SV_T �  $CUR_SV_ANG   	��ARMLOAD_T �  $ARMLOAD   t�ARMLOAD_P_T �  $ARMLOAD_P    H�MRR2_GRP_T �� $ARM_PARAM   d$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$RLIBSW01  $RLIBSW02  $ABC_FLAG  $MD_J2SECT   $MD_J3SECT   
$MD_J1SPCONS   P$MD_J2SPCONS   P$MD_J3SPCONS   P$MD_CUR_K   $MD_CUR_J2  $MD_CUR_J3  $SV_OFF_TIM2   	$CSKPLIM_ENB  $CSKPLIM_LIN  $CSKPLIM_JNT   	$QSKPLIM_ENB  $QSKPLIM_LIN  $QSKPLIM_JNT   	$EXT_AZIM   $EXT_ELEV   $SERVOCMPTOL   	$ARMLOAD 1� $ARMLOAD_X 1� $ARMLOAD_Y 1� $ARMLOAD_Z 1� 	��INTERACT_T �  $INTERACTION   	�INTRAC_N_T �  $INTRAC_NUM   	��INTRAC_D_T �  $INTRAC_DIV   	��DH_EXTRA_T � 0 $VALID  $X  $Y  $Z  $W  $P  $R  �MRR_GRP_T �H �$BELT_ENABLE  $CART_ACCEL1  $CART_ACCEL2  $CIRC_RATE  $CONTAXISNUM  $PS_EXP_ENBL   $EXP_ENBL  $JOINT_RATE  $LINEAR_RATE  $PATH_ACCEL1  $PATH_ACCEL2  $PATH_ACCEL3   $PROCESS_SPD  $PROC_SPDLIM  $CNT_ACC_MGN  $DDACC_RATIO  $FWP_TIME1  $FWP_TIME2  $ACCEL_RATIO  $DECEL_RATIO  $PPABN_ENBL  $ROTSPEEDLIM  $SPEEDLIM  $SPEEDLIMJNT  $DEF_MAXACCE   $USE_CAL  $SPIN_CTRL  $SYN_ERR_LIM   $SYNC_GAIN   $SYNC_OFFSET   $MOUNT_ANGLE  $COLLINEAR  $COINCIDENT  $ACCEL_TIME1   	$ACCEL_TIME2   	$ENCSCALES   	$EXP_ACCEL   	$PS_INPOS_TI   $INPOS_TIME   	$JNTVELLIM   	$JNT23_UPLIM  $JNT23_LOWLI  $LOWERLIMS   	$LOWERLIMSDF   	$MASTER_POS   	$MIN_ACCTIME   	$MOSIGN   	$MOT_SPD_LIM   	$PERCH    	$MOVERRLIM    	$PERCHTOL    	$STOPERLIM   	$STOPTOL   	$SERVO_CTRL  $PS_SV_OFF_A   $SV_OFF_ALL  $SV_OFF_ENB   	$SV_OFF_TIME   	$UPPERLIMS   	$UPPERLIMSDF   	$TRKERRLIM  $PAYLOAD  $PS_MAX_PAYL   $MAX_PAYLOAD  $AXISINERTIA   	$AXISMOMENT   	$MAX_AMP_CUR   	$ACCEL_PARAM   $MAX_PTH_ACC  $MRRDUM2   $PS_BCKLSH_C   $BCKLSH_COUN   	$MOVER_GAIN   	$MOVER_SCALE   	$MOVER_OFFST   	$CLALM_TIME  $TSMOD_TIME  $CHKLIMTYP  $SNGLRTY_STP  $INPOS_TYPE  $JOG_TIME_M  $MIN_ACC_UMA  $MIN_ACC_UCA  $ACC_SCL_UCA  $SLMT_J1_LW   $SLMT_J1_UP   $SLMT_E1_LW   $SLMT_E1_UP   $SLMT_J1_NUM  $SLMT_E1_NUM  $PS_SPCCOUNT   $SPCCOUNTTOL   	$SPCMOVETOL   	$SHORTMO_MGN  $MIN_ACC_CMC  $EXTACCRATIO  $CN_GEAR_N1  $CN_GEAR_N2  $SFLT_ERLIM   	$SV_CTRL_TYP   	$PS_CARTMO_M   $CARTMO_MGN  $MIN_CAT_UMA  $MIN_ACC_SHM  $GEAR_RATIO   	$EXP_JOG_ACC   	$PS_ARMLOAD   $ARMLOAD   $ACC_PA_UMA  $ACC_PC_UMA  $AXIS_IM_SCL  $PS_MOT_LIM_   $MOT_LIM_STP  $JG_FLTR_SCL  $JOGACCRATIO   $TORQUE_CONS   	$MIN_PAYLOAD  $DECOUP_MGN   $DECP_MGN_WR   	$PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $FFG_MGN_J2  $FFG_MGN_J3  $DVC_AC0_MAX   	$DVC_AC1_MAX   	$DVC_ACC_MAX   	$DVC_ACC_MIN   	$DVC_JRK_MAX   	$DVC_JRK_MIN   	$SV_DBL_SMT  $SV_MCMD_DLY  $SV_GRV_X  $SV_GRV_Y  $SV_GRV_Z  $SV_DH_D   	$SV_DH_A   	$SV_DH_COSA   	$SV_DH_SINA   	$SV_LNK_M   	$SV_LNK_X   	$SV_LNK_Y   	$SV_LNK_Z   	$SV_LNK_IX   	$SV_LNK_IY   	$SV_LNK_IZ   	$SV_Z_SIGN   	$SV_DMY_LNK   	$SV_DH_COSTH   	$SV_DH_SINTH   	$SV_THET0   	$LNK23Z  $LNK23X  $LNKCBZ  $LNKCBX  $CB_MASS  $CB_IX  $CB_IY  $CB_IZ  $LNKSBY  $LNKSBX  $LNGTSB  $SPCNS  $ARMLOAD_X   $ARMLOAD_Y   $ARMLOAD_Z   $DUTY_ENB   	$DUTY_PARAM1   	$DUTY_PARAM2   	$QSTOP_TOL   	$NE_ENB  $LINK_TYPE   	$ARMLOAD_NUM   	$DH_THETA0   	$DH_THETA   	$DH_D   	$DH_A   	$DH_ALPHA   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	$DH_VD   	$DH_VA   	$DH_VALPHA   	$LINK_VM   	$LINK_VSX   	$LINK_VSY   	$LINK_VSZ   	$LINK_VIX   	$LINK_VIY   	$LINK_VIZ   	$DH_HD   	$DH_HA   	$DH_HALPHA   	$LINK_HM   	$LINK_HSX   	$LINK_HSY   	$LINK_HSZ   	$LINK_HIX   	$LINK_HIY   	$LINK_HIZ   	$DH_OTHETA   	$DH_OD   	$DH_OA   	$DH_OALPHA   	$LINK_OM   	$LINK_OSX   	$LINK_OSY   	$LINK_OSZ   	$LINK_OIX   	$LINK_OIY   	$LINK_OIZ   	$FLINK_BX   	$FLINK_BY   	$FLINK_BETA   	$SPBALANCE_K   	$SPLENGTH_0   	$SPACT_X   	$SPACT_Y   	$SPACT_Z   	$SPFULC_X   	$SPFULC_Y   	$SPFULC_Z   	$INTERACTION 1� 	$AUTO_SNGSTP  $T1T2_SNGSTP  $CART_2ND_TI  $JNT_2ND_TIM   	$LC_QSTP_ENB  $CP_CUTOFFOV  $CP_MINSEG  $MASTREV_ENB  $MASPOS_DIFF   	$INTRAC_NUM 1� 	$INTRAC_DIV 1� 	$OBS_DIST  $SV_PARAM   2$MIJNTCHKLMT  $LCHWARN_ENB  $ABC_PARAM   $MECH_MASK  $MECH_TYPE  $AXS_MAP_NUM  $AXS_MAP   	$DH_EXTRA 1� 
$AXS_COUPLE   	$PS_ROBOT_CR   $ROBOT_CRC  �0�MSK_CE_GRP_T � P $T1_USERCART  $T1_USERJNT   	$T1_CARTVEL  $T1_JNTVEL   	$T1_WARNING  �MTCOM_CFG_T �  $CNC_NO  $NORES_TIMEO  �OPWORK_T �, $SYSBUSY  $SOPBUSYMSK  $TPBUSYMSK  $UOPBUSYMSK  $INTPRUNNING  $INTPPAUSED  $INTPMASK  $OPT_OUT  $UOP_DISABLE  $OUTIMAGE   $OP_PREV_IMG   $OP_INV_MASK   $ORGOVRDVAL  $USER_OUTPUT   $PS_ENBL_ON   $ENBL_ON  $MLT_RBT_ENB  $PMC_EDT_MSK   $NOALM_MSK  $DUMMY19  ! �OVRDSLCT_T � x $OVSL_ENB  $SDI_INDEX1  $SDI_INDEX2  $OFF_OFF_OVR  $OFF_ON_OVRD  $ON_OFF_OVRD  $ON_ON_OVRD  $DUMMY   5��OVRD_SETUP_T � @ $OVRD_NUM  $OVERRIDE   
$OVRD_NUM_S  $OVERRIDE_S   
 ��TRACECTL_T � H $TASK_STATUS  $TRC_TOP_IDX  $TRC_BTM_IDX  $TASK_ID  $DUMMY4  �TRACEDT_T � D $EPT_INDEX  $LINE_NUM  $FILE_OFST  $EXEC_TYPE  $LINE_ST  �TRACEUP_T � @ $TRC_UPDATE  $DISP_PXNN  $DUMMY2  $DUMMY3  $DUMMY4  ��PG_CFG_T � $SUBTASKNUM  $NUM_TASKS  $JMPWAIT_UPR  $JMPWAIT_LOW  $FAST_MODE  $RCVFAIL_CNT  $WAITREL_CFG  $ACC_CTRL  $CNT_CTRL  $IGNR_PLS  $DBTB_STPTYP  $BWD_CFG  $RESUME_CFG  $IGPAUS_PRI  $MTNLN_CFG  $PAUS_RTN  $RESERVE1  $RESERVE2  ��PG_DEFSPD_T � L $AP_DEF_SPD  $AP_DEF_UNIT  $DUMMY4  $APSP_PREXE  $DLY_LASTPS   ��PING_T � 0 $TIMEOUT  $DATALEN  $NPACKETS  $DEBUG  �PIPE_CFG_T � h $ARSIZE   $FILEDATA   $SECTORS  $FORMATTER  $RECORDSIZE  $MEMTYPE  $FORMAT  $AUXWORD   	��PLID_CFG_T �  $COMP_SWITCH   T�MAX_PLD_CAL_ � $ $AA  $BB  $CC  $DD  $EE  �CALC_RESULT_ � � $PAYLOAD  $PLD_J3ARM  $INERTIA4  $INERTIA5  $INERTIA6  $MOMENT4  $MOMENT5  $MOMENT6  $COMB_LOAD4  $COMB_LOAD5  $COMB_LOAD6  $PUB_INRT4  $PUB_INRT5  $PUB_INRT6   P�PLID_GRP_T �P H$PI_ENB  $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $ARMLOAD3  $ROB_TYPE  $DATA_NUM  $SPEED_HIGH  $SPEED_LOW  $DEFSPD_HIGH  $DEFSPD_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DEFACC_HIGH  $DEFACC_LOW  $SAMPLE_TIME  $SAMPLE_HIGH  $SAMPLE_LOW  $MOV_AXIS   	$MOV_POS1   	$MOV_POS2   	$MOV_DEF1   	$MOV_DEF2   	$ROT_INERTIA   	$MAX_VEL_HI   	$MIN_VEL_HI   	$MAX_ACC_HI   	$MIN_ACC_HI   	$MAX_VEL_LOW   	$MIN_VEL_LOW   	$MAX_ACC_LOW   	$MIN_ACC_LOW   	$GAMMA   	$STOP_DATA  $GETDATA_FIN  $ID_RESULT   
$CALIBRATE  $PI_DEBUG  $HIDAT_V_MAX   	$HIDAT_V_MEA   	$HIDAT_A_MAX   	$HIDAT_A_MEA   	$LWDAT_V_MAX   	$LWDAT_V_MEA   	$LWDAT_A_MAX   	$LWDAT_A_MEA   	$CALC_TYPE  $MTN_CALCTYP  $CHKER_VER $PDCK_RB_TYP  $I_FACTOR   $MAX_PAYLOAD  $MAX_INERTIA   $MAX_MOMENT   $COMB_LOAD   $MAX_PLD_CAL �$IM_SRCH_DT  $WARN_DISP  $WARN_LEVEL  $OVER_LEVEL  $CALC_RESULT �$PAMSWFLG  $AMLD_SCRN  $DUMMY69  $DUMMY70  $DUMMY71   ��PLID_SV_T �P $CUR_SCRN  $CUR_GROUP  $PS_SAVE_DON   $SAVE_DONE  $NO_RECOVER  $RESULT_SAV   
$PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $DO_DEFAULT  $MOV_POS1   	$MOV_POS2   	$SPEED_HIGH  $SPEED_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DO_DEF_POS   `�PLIM_GRP_T � � $MAX_PYLD  $AXISINERTIA   	$AXISMOMENT   	$AXIS_IM_SCL  $PS_LIM_WT_S   $LIM_WT_SCL  $LIM_INR_SCL   $LIM_MNT_SCL   $LIM_CL_SCL   $PLD_MODE  $DUMMY10  $DUMMY11  h�PLMR_GRP_T � � $PYLD_ENB  $WMR_ENB  $ANGLE  $PLMR_AA  $PLMR_BB  $PLMR_CC  $PLMR_DD  $PLST_ANG   
$COMP_SW  $MAX_XY_LOC  $MAX_Z_LOC  �PLST_GRP_T � p $COMMENT $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  �PL_RES_G_T � | $PAYLOAD  $SAVMOMENT4  $SAVMOMENT5  $SAVMOMENT6  $SAVINERTIA4  $SAVINERTIA5  $SAVINERTIA6  $EST_RESULT   0��PL_RES_V_T �  $PL_RES_G_P   �PMON_QUE_T � 8 $QCOUNT  $QTHRESHOLD  $QHYSTERESIS  $QUEUE_UP  �PM_GRP_T � � $ACC_TIME1  $ACC_TIME2  $POS_ERR_LIM  $ROT_ERR_LIM  $ENABLED  $DBG_MASK  $COMP_SWITCH  $BWD_ACC1  $BWD_ACC2  $JVEL_RATIO  $REWIND_NUM  $GTF_ACC1  $GTF_ACC2  �POCFG_T �   $PODEBUG  $OVERRUN_TOL   �PODATA_T � P $OVERRUN_CNT  $CUR_INDEX  $PROGRAM_ID   2$LINE_NO   2$OVERRUN_ITP   2�POINFO_T �  $CUR_INDEX  $INFO   ���POIO_T � ( $SLEQ_NUM  $IO_TYPE  $IO_INDEX  ��POS_EDIT_T � � 	$LOCK_POSNUM  $HIDE_MENU  $HIDE_POSNUM  $AUTO_RENUM  $COPY_POSDAT  $AUTO_RENUM2  $RMV_MANRENM  $COPY_POSTYP  $CPRUT_ENB   �PRGADJ_T � h $X_LIMIT  $Y_LIMIT  $Z_LIMIT  $W_LIMIT  $P_LIMIT  $R_LIMIT  $SPEED_ADJ  $NEXT_CYCLE  ��PRGNS_CFG_T � � $ALGO_VER  $NYQ_FREQ  $WIN_TYPE  $WIN_SIZE  $OVERLAP  $FREQ_LIM  $MIN_NUM  $CREATED  $VERIFY  $PROGNAME %$CREATE_GP  $STATUS_GP  $DEBUG  $MAILTIME  $MAILEVENT  $LASTMAIL  �PRGNS_ELEM_T � � $ENABLE  $FEASIBLE  $AXIS  $PS_ELEM_NUM   $ELEM_NUM  $ROT_RATIO  $MAX_FREQ  $THRE_REL  $THRE_ABS  $DEGRAD_LVL  $DEGRAD_BASE  $DEGRAD_RATE  $UPD_DATE $BASE_DATE P��PRGNS_GRP_T � X $ELEM 2� $MIN_ANG   	$MAX_ANG   	$BASE_ANG   	$LAST_MOD   	$BASE_MOD   	 
��PRGNS_PREF_T � ( $GRIDLINES  $BARS_NUM  $STYLE  ��PROTOENT_T �  $P_NAME !$P_PROTO  �PROXY_CFG_T � � $LIST_PORT  $PROXY_ENB  $PROXY_SRV )$PROXY_PORT  $DIRECT_1 )$DIRECT_2 )$DIRECT_3 )$DIRECT_4 )$DIRECT_5 )$DIRECT_6 )$DIRECT_7 )$DIRECT_8 )T�PF_DATA_T �   $VALUE  $GROUP  $AXIS  
��PF_CFG_T �| $ENABLE  $PROG_NAME %$CUR_GROUP  $RAN_GROUPS  $START_TYPE  $TOTAL_TIME  $TOTAL_PWR  $INS_PWR  $REGEN_PWR  $INS_REGEN  $EXE_DATE $DATA_TYPE  $RES_NAME %$MONTR_RATE  $D_PWR_SUP  $D_PWR_REG  $RV_LIM1  $RV_LIM2  $DEGREE  $REFRESH  $OVERRIDE  $RV_HRS_DAY  $RV_DAYS_YR  $MAXSIZE  $SUMMARY 2� $CONFIG_SET  $SUPPORT  $LAST_RUN   ,�PF_PREF_T � 4 $GRIDLINES  $BARS_NUM  $DATA_TYPE  $STYLE  �PSSAVE_T � $MC_FOLDER 	$SLAVE_SAVE  $START_MULTI  $SLAVE_LOAD   $LOAD_DEV  $KEEP_HNADDR !$KEEP_HRADDR !$KEEP_CCOMM $KEEP_CPROT 	$PS_KEEP_COP   $KEEP_COPER  $KEEP_CSTATE  $KEEP_CREMOT $KEEP_CTIMEO  $KEEP_CSREMO $KEEP_CUNAME e$KEEP_CHPWD  $KEEP_SBMSK !d�PSSAVE_GRP_T � , $FLANGE  $SYNC_FLANGE  $SYNC_MST_CN  �PS_CONFIG_T � � $DB_IMMTRIG  $DA_IMMTRIG  $DB_NOTRIG  $DA_NOTRIG  $TCLAMP_WARN  $USE_DYNSPD  $MAX_SEARCH  $NUM_PSMOTN  $DB_MARGIN  $RESOLUTION  $COMP_MASK  $PX_STARTED  $SCAN_READY  $SCAN_ALIVE  �PS_CP_CFG_T �  $ENB  $REF_MODE  ��PS_CP_GRP_T � � 
$ENB  $REF_MODE  $FLANG_VALID  $FLANG_TICK  $FLANG_TRANS $PREVI_TRANS $UTOOL_VALID  $UTOOL_TRANS $FKSOL_FP  $SEG_COUNTER   �PS_ITEM_T � � $BASE_DIST  $TUNE_MSEC  $MN_LEN  $ITEM_LINE  $ITEM_DONE  $TRIGGERED  $STOP_TRIG  $NG_ITEM  $CLAMPED  $PARAM1  $PARAM2  $PARAM3  $ML_ACT_P  $MN_CODE   �PS_MOTION_T ��  $OWNER_TID  $G0  $PS_DONE  $PG_STATUS  $DB_STATUS  $DA_STATUS  $DB_MIN_DIST  $DA_MAX_DIST  $PARENT_NAME %$CHILD_NAME %$PARENT_LINE  $SCAN_COUNT  $SEG_STARTED  $SEG_COUNTER  $SCAN_ABORT  $PARENT_EPT  $CHILD_EPT  $PRV_VALID  $PRV_DB_DIST  $PRV_DA_DIST  $PRV_VEC   $PRV_TICK  $BASE_SPEED  $DEST_VALID  $DEST_VEC   $UT_TRANS $MMR_P  $MODONE  $NEXT_MODONE  $SMH_MASK  $NUM_ITEM  $ITEM 2� ��PWRUP_DLY_T �   $DELAY_TIME  $SY_READY   
��QSKIP_GRP_T � � $ERROR_CNT2   	$QSKP_ERRCNT   	$QSKP_CURANG  $QSKP_CURAN1  $QSKP_CURAN2  $QSKP_CURAN3  $QSKP_CURAN4  $QSKP_CURAN5  $QSKP_CURAN6  $QSKP_CURAN7  $QSKP_CURAN8  $QSKP_CURAN9  �J2RED_T � 4 $EXD_RTQ  $EXD_ITP  $EXD_PRG  $EXD_LINE   (�RDCR_GRP_T � � $RMAX_TORQUE   	$RMIN_TORQUE   	$THRES_TORQ   	$RGEAR_RATIO   	$WARN_FLG   $COMP_SW  $RESERVE   	$SPC_ITP  $NUM_EXD  $J2TH2ND  $J2RED 1� ��REFPOS11_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS21_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS31_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS41_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS51_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS61_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS71_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS81_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPSMSK_T �  $MAXREFPOSEN    ��REMOTE_CFG_T � 4 $REMOTE_TYPE  $REMOTEIOTYP  $REMOTEIOIDX   `�REPOWER_T �  $FLAG  ��RESTART_T � , $FLAG  $DSB_SIGNAL  $STARTUP_CND   ��RS232_CFG_T � � $COMMENT $DEVICEUSE  $SPEED  $PARITY  $STOPBITS  $FLOWCONTROL  $TIMEOUT  $CUSTOM  $AUXTASK  $INTERFACE  $STATUS  ��RSCH_T � @ $OLD_SPEC_SW  $FREEFROMSIZ  $TARGET_DIR 	$UPDT_MAP   L�RSPACE_T �� !$COMMENT $USAGE  $ENABLED  $IN_EXTERIOR  $ENTRY  $ENT_SIGN_ON  $PRIORITY  $PRIORWRK  $DOUT_TYPE  $DOUT_INDX  $DIN_TYPE  $DIN_INDX  $FRIEND_GRP  $UFRAM_NUM  $UTOOL_NUM  $MYHOLD  $LENGTH_VTEX  $FIRST_VTEX   $SECND_VTEX   $UFINV_POST $MARGIN  $WAITING  $FIRST_VTX2   $SECND_VTX2   $G2ENTRY  $G1ENT_INTR  $G2ENT_INTR  $PRE_UFRAM  $NO_USE_DI  $HOLD_REQ  $CSPACE_NUM  $CUR_TCP   $PRE_TCP   h�GP_STATUS_T � @ $IN_USE  $SPACE_NUM  $PRIORITY  $STATUS1  $STATUS2  \�COM_SPACE_T �X $USE_MLT_CTN  $H_PRIORITY  $IN_CONTROL  $IN_SPACE_GP  $WT_SPACE_GP  $USE_GP  $DEADLOCK_GP  $DELAY_CNT1  $DELAY_CNT2  $GP_STATUS 2� $DOUT1_TYPE  $DOUT1_INDX  $DOUT2_TYPE  $DOUT2_INDX  $DOUT3_TYPE  $DOUT3_INDX  $DIN1_TYPE  $DIN1_INDX  $DIN2_TYPE  $DIN2_INDX  $EXT1  $EXT2  $V1   $V2   $V3   ��GP_HOLD_T � � $STATUS  $GP_MSK  $SPACE_NUM  $CSPACE_NUM  $REQ_GRP  $PS_RATE   $RATE   $INT_POS   $ACT_POS   $PRD_POS   $S1  $S2  $S3  $S4   x�RSPACEG_T � 0 $COM_SPACE 2� $GP_HOLD 2� $SPARE_INT   
 �RSPACESR_T � � $SR_ENB_TYP   $RUNNER_AXS  $HAND_LNGTH  $HAND_THICK  $FLIP_ENB  $INTFERENCE  $HAND_IF_CHK  $HANDI_TYPE  $HANDI_INDX  $SR_G1POS   $SR_G1POS_IN   $SR_G1ANG   $SR_G1ANG_JF   $SR_PRM   	�RTCFG_T � � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $RSM_RTCP  $INLINE_WRST   $TBC_PTH_CMP  $DRTCP_ENB  $LDR_SP_RATE  $LDR_RSP_RAT  $COMP_SWITCH   8�RV_DATA_T �  $DATETIME    	$VALUE    	�RV_DATA_GRP_ �  $DATA  2� �SCR_T �	| �$ITP_TIME  $NUM_GROUP  $NUM_TOT_AXS  $NUM_DSP_AXS  $JOGLIM  $FINE_PCNT  $COND_TIME  $MAXNUMTASK  $KEPT_MIRLIM  $MAXPREMTN  $MAXPREAPL  $PRE_EXE_ENB  $NUM_SYS_MIR  $NUM_PG_MIR  $BRKHOLD_ENB  $ENC_AXIS    $ENC_TYPE    $NUM_GP_MADE  $NUM_RLIBSOC  $NUM_MOTNSOC  $DUMMY158  $SV_CODE_OPT  $SFSPD_OVRD   $COLDOVRD  $COORDOVRD  $TPENBLEOVRD  $FENCEOVRD  $JOGOVLIM  $SFJOGOVLIM  $RUNOVLIM  $SFRUNOVLIM  $MAXNUMUFRAM  $MAXNUMUTOOL  $LCHDLY_TIME  $RECOV_OVRD  $JOGWST_MODE  $JOGLIMROT  $MOTN_PC_RUN   @$RESETINVERT  $OFSTINCVAL  $FWDENBLOVRD  $TPMOTNENABL  $PREV_CTRL  $MAX_PRE_FDO  $PRE_MB_CMP  $MB_DSBL_MSK  $MB_DSB_MSK2  $SVSTAT  $UPDATE_TIME  $JG_DSBL_MSK  $NUM_PG_AMR  $MB_LD_MSK  $MOTN_LD_MSK  $MOTN_LD_MK2  $AMP_TYPE   T$CAP_AMP_DIS   T$HBK_MAP_ENB  $HBK_IO_TYPE  $HBK_IO_IDX  $PPA_MAP_ENB  $PPA_IO_TYPE  $PPA_IO_IDX  $MOTN_LD_IDX   @$DVC_DBG  $DVC_ENB  $DVC_MODE  $DVC_MODE1  $DVC_MODE2  $DVC_MODE3  $DVC_C_RATIO  $INTASK_OVRU  $DSP_TYPE  $CABINET_TYP  $NE_MODE  $PG_DSBL_MSK  $JOG_AUX_ENB  $SUBCPU  $NE_SIN_RESO  $UPDATE_MAP1  $UPDATE_MAP2  $UPDATE_FLAG   $HW_C1_TIME1  $HW_C1_TIME2  $ATR   �$UNITTYPE   �$ATRATTRIB   �$NE_CYCLE  $NECA_OVRUN  $FLTR_2_FIX  $STARTUP_CND  $DSB_SIGNAL  $LPCOND_TIME  $CHK_CH_SCTM  $F_ATR   �$F_UNITTYPE   �$F_ATRATTRIB   �$FSSB_STAT   �$CHAIN_TIME  $CHAIN_STAT  $CHAIN_RSDN  $DSP_MAP_ENB  $IDX_TBL_MSK  $PROC_CTRL  $TEMPER_LIMS   T$FSSB1   $FSSB2   $FSSBDIAGENB  $RAILACC_ENB  $SMCR_LOADED  $DUMMY159  $PS_DSP_TYPE   $DSP_TYPE2  $PRC_DSP   $PRC_CD_ID 	$MOTN_FUNC   $INTRINS_TP  $DIAG_FUNC  $TRANS_NUM   T$TRANS_MAX   T$TRANS_WARN   T$CBLCUR_MAX   T$CBLCUR_A   T$CBLCUR_B   T$CBLCUR_WARN   T$DAC_TRANS   T$DAC_CBLCUR   T$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $CE_RIA_SW  $SAFE_SPD  $SAFE_ROTSPD  $T2_LOCK_ENB  $DSB_MOINIT  $MAX_DF_LEN  $MPDT_TIMLMT  $FAST_HRDYON  $ORG_PTH_RSM  $DAC_LMT  $MULSELENB  $UPDATE_MAP3   $JCOLDOVRD  $JTPENBOVRD  $JFENCEOVRD  $FAN_ALMLVL  $FAN_WRNLVL  $HARDTYP_MAP  $COMP_SW   2$SHADOWRECS  $SHADOWTIME  $FANSTOP_TIM  $BRK_ECO_ENB  $AUTATR_STAT  $AUTO_SBRIDX  $AUTO_DSPIDX  $AUTO_ATRIDX   $AUTO_AMPINF   �$AUTO_AMPCUR   �$REGTYPE  �AX_OFS_T �  $X  $Y  $Z  <�SCR_GRP_T �� �$NUM_SEG   $NUM_PT   $ARM_TYPE  $DUMMY121  $ARM_TYPE_B  $NUM_AXES  $NUM_ROB_AXS  $NUM_RED_AXS  $WRST_AXIS_S  $WRST_AXIS_E  $SYNC_M_AXIS  $SYNC_S_AXIS  $WRIST_TYPE  $HW_STRT_AXS  $AXISORDER   	$DUMMY122  $BRK_NUMBER   	$DUMMY123  $DD_MOTOR   	$ROTARY_AXS   	$LOADRATIO   	$CONFIG_MASK  $LINK_LENGTH   $EXT_ORDER   $DUMMY124  $EXT_XYZ_MAP   $DUMMY125  $EXT_OFFSET   $EXT_LENGTH   $ROBOT_ID $ROBOT_MODEL 	$ROBOT_FILE 	$ROBOT_INT  $SV_CODE_ID $JOGLIM_JNT   	$COORD_MASK  $OP_BRK_NUM   	$DUMMY126  $USE_TBJNT  $USE_TBCART  $NUM_DUAL  $DUMMY127  $PS_TURN_AXI   $TURN_AXIS   $AXS_AMP_NUM   	$FLEXTOOLTYP  $AXS_XYZ_MAP   	$DUMMY128  $OFST 1� 	$KINEM_ENB  $DUMMY129  $PS_UPDATE_M   $UPDATE_MAP  $TORQCTRL  $DSP_NUM   	$DUMMY130  $PS_M_POS_EN   $M_POS_ENB  $M_DST_ENB  $MOVE_DST  $MCH_POS_X  $MCH_POS_Y  $MCH_POS_Z  $MCH_POS_W  $MCH_POS_P  $MCH_POS_R  $MCH_ANG   	$MCH_SPD  $DST_MIR_P  $DPOS_DST  $DST_POS_X  $DST_POS_Y  $DST_POS_Z  $DSP_ERCNT   	$PS_DEST_DAT   $DEST_DATA_P   $ROBOT_FUNC  $PROC_AXS   	$DAC_MODE  $DAC_AXMODE   	$DAC_RATE1   	$DAC_RATE2   	$DAC_RATE3   	$DAC_RATE4   	$DAC_RATE5   	$DAC_RATE6   	$DAC_RATE7   	$DAC_RATE8   	$DAC_RATE9   	$DAC_RATE10   	$DAC_LMT1   	$DAC_LMT2   	$DAC_LMT3   	$DAC_LMT4   	$DAC_LMT5   	$DAC_LMT6   	$DAC_LMT7   	$DAC_LMT8   	$DAC_LMT9   	$DAC_LMT10   	$DAC_DEBUG   $FUNC_SW   $FUNC_VAL   $ABC_ENB  $HBK_ENBL  $MV_DIAG   
$ABC_MODE1  $ABC_MODE2  $ABC_MODE3  $ABC_MODE4  $ABC_MODE5  $ABC_MODE6  $ABC_MODE7  $ABC_MODE8  $ABC_MODE9  $SAFE_JNTSPD   	$ROBOT_LABEL $DSP_NUM_FLG  $GROUP_NUM  $COMP_SW   $AMB_TEMP  $DSP_STRT_AX  $TOT_SBR_NUM  $TOT_DSP_NUM  $TOT_ATR_NUM  $TANDEM_SUB   	$DSP_ORDER   	$ATR_ORDER    $AMPINF_ORDR    $AMPCUR_ORDR    $FIX_ORNT_WR  �SERVENT_T � $ $S_NAME !$S_PORT  $S_PROTO !��SERV_MRA_T � d $DATETIME  $ERR_CODE  $SAFETY_ST  $IMP_VEL   	$IMP_TOQ   	$ANGLES   	$DIST_TOQ   	 ��SERV_REC_GRP � p $TOTAL  $BIN_V1T1   	$BIN_V1T2   	$BIN_V2T1   	$BIN_V2T2   	$MRA_REC 1� 
$MRA_IDX  $WCA_REC 1� 
��SERV_RV_T �  $OVER_LIMIT   	��SERV_OCCUR_T �  $ERR_CODE  $COUNTER   �SHELL_CFG_T � 5$JOB_BASE  $RSR_ENABLE   $NUM_RSR   $RSR1_NAME %$RSR2_NAME %$RSR3_NAME %$RSR4_NAME %$RSR5_NAME %$RSR6_NAME %$RSR7_NAME %$RSR8_NAME %$JOB_ROOT %$CONT_ONLY  $USE_ABORT  $RSR_ACKENBL  $INVERT_CHK  $UOP_SEL_STA  $RSR_ACK_PUL  $COM_TIMEOUT  $PNS_ENABLE  $SHELL_NAME %$START_MODE  $TPFWD_KAREL  $ERR_REPORT  $OPTIONS  $QUE_ENABLE  $PRODSTARTYP  $CSTOPI_ALL  $SHELL_EXT  $SEL_TYPE  $EXT_SEM1  $EXT_SEM2  $MAINT_STYL  $ISOL_ENB  $DI_CHKTRIG  $PROD_MODE  $INIT_TMO  $MANRQ_TMO  $EXTEND_ENB  $KEYSWITCH  $STARTCHKTYP  $HEARTBEATMS  $PERM_LEVEL  $TEMP_LEVEL  $USTART_FT  $START_SIG  $DO_HOME_SOP  $REFPS_PR_ID  $DIS_STRTCHK  $CUSTOM  $E_RECOV_MSK  $SET_IOCMNT  $CSTOPI_ALL2   \�SHELL_CHK_T � D $ENABLE  $RESUME  $PROMPT  $ERRPOST  $FORCE  $WARN   ��SHELL_COMM_T � @ $FUNC  $STATUS  $PARM1  $PARM2  $PARM3  $PARM4   ��SMB_HDDN_T �  $BLOB    �SNPX_ASG_T � 0 $ADDRESS  $SIZE  $VAR_NAME %$MULTIPLY  �SNPX_PARAM_T � � $TIMEOUT  $SNP_ID 	$NUM_ASG  $NUM_CIMP  $NUM_FRIF  $VERSION  $STATUS  $DISP_INFO  $MODBUS_ADR  $NUM_MODBUS  $MODBUS_PORT   ��SSR_T � x $SINGLESTEP  $DUMMY7  $SGLSTEPTASK   &$STEPTASKNUM  $STEPSTMTTYP  $STPSEGTYPE  $BWDSTEP  $SHOWSTMTTYP  �SVDT_GRP_T �� �$DATA00   	$DATA01   	$DATA02   	$DATA03   	$DATA04   	$DATA05   	$DATA06   	$DATA07   	$DATA08   	$DATA09   	$DATA0A   	$DATA0B   	$DATA0C   	$DATA0D   	$DATA0E   	$DATA0F   	$DATA10   	$DATA11   	$DATA12   	$DATA13   	$DATA14   	$DATA15   	$DATA16   	$DATA17   	$DATA18   	$DATA19   	$DATA1A   	$DATA1B   	$DATA1C   	$DATA1D   	$DATA1E   	$DATA1F   	$DATA20   	$DATA21   	$DATA22   	$DATA23   	$DATA24   	$DATA25   	$DATA26   	$DATA27   	$DATA28   	$DATA29   	$DATA2A   	$DATA2B   	$DATA2C   	$DATA2D   	$DATA2E   	$DATA2F   	$DATA30   	$DATA31   	$DATA32   	$DATA33   	$DATA34   	$DATA35   	$DATA36   	$DATA37   	$DATA38   	$DATA39   	$DATA3A   	$DATA3B   	$DATA3C   	$DATA3D   	$DATA3E   	$DATA3F   	$DATA40   	$DATA41   	$DATA42   	$DATA43   	$DATA44   	$DATA45   	$DATA46   	$DATA47   	$DATA48   	$DATA49   	$DATA4A   	$DATA4B   	$DATA4C   	$DATA4D   	$DATA4E   	$DATA4F   	$DATA50   	$DATA51   	$DATA52   	$DATA53   	$DATA54   	$DATA55   	$DATA56   	$DATA57   	$DATA58   	$DATA59   	$DATA5A   	$DATA5B   	$DATA5C   	$DATA5D   	$DATA5E   	$DATA5F   	$DATA60   	$DATA61   	$DATA62   	$DATA63   	$DATA64   	$DATA65   	$DATA66   	$DATA67   	$DATA68   	$DATA69   	$DATA6A   	$DATA6B   	$DATA6C   	$DATA6D   	$DATA6E   	$DATA6F   	$DATA70   	$DATA71   	$DATA72   	$DATA73   	$DATA74   	$DATA75   	$DATA76   	$DATA77   	$DATA78   	$DATA79   	$DATA7A   	$DATA7B   	$DATA7C   	$DATA7D   	$DATA7E   	$DATA7F   	 4�SVPRM_UPD_T �  $PRM   
��SVGUN_CT_T � ` $OUTPUT_ENB  $INPUT_ENB  $GROUP_NUM  $AXIS_NUM  $GO_VALUE  $GI_VALUE  $IO_SCALE  �SYSLOG_T � � $SIZE  $MODE  $STATUS  $ADDRESS  $DATA_SIZE  $COMP_VALUE  $STOP_MODE  $CURR_VALUE  $FLOG_ID_LO  $FLOG_ID_HI  $FLOG_ID_IN  $FILE_OUT  $FILE_NAME $ID  ��SYSLOG_SAV_T � h $SAVE_BLCKS  $SAVE_TASKS  $SAVE_D_CPU  $SAVE_D_SIZ  $SAVE_D_ADD  $FILE_OUT  $FILE_NAME �SYSTEM_TIMER � p 
PWR_TOT  PWR_LAP  SRV_TOT  SRV_LAP  RUN_FLG  RUN_TOT  RUN_LAP  WIT_FLG  WIT_TOT  WIT_LAP  �TBC_ACC_T �X -$ACC_LEN1  $ACC_LEN2  $ACCEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT   	$M_STAT  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $AC_ACC  $JK_ACC  $VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AAL1  $AAL2  $AAL3  $AAL4  $AAL5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM   2$�TBCCFG_T � ` $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $TBC_STAT   $TC 2� $TBC_DEBUG  �TBCSG_GRP_T � \ $ENABLE  $APPRC_SCL   
$OPEN_SCL   
$CLOSE_SCL   
$CLS_MINF2   
$CLS_MINACC   
�$$CLASS  ������       �$$VERSION  ������  ���$AAVM_WRK 2 ������ 0  �5�                                �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            T  �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                              �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            AC_D�                                                 	 	                                     ���� 	                                     ����                                                       	                                                             �$ABSPOS_GRP 1������� <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �$ACC_MAXLMT         ��   ��$ACC_MINLMT        ��    �$ACC_PRE_EXE        ��    �$AC_UPDATE  �����������$ALARMRECOV ������   �        �$ALMDG ������                �$ALM_IF ������    d                                                                                                       d                                                                                                         , 
                                         �$ANGTOL  ������� 	 A   A   A   A   A   A   A   A   A   �$APPLICATION ?������� 
 HandlingTool          
V8.20P/A2          �� 
88150              ���
3347126            �  
471                ���
V8.20P/A2             7DE3/A2               	80604.015             FRL                ���2                   �$AP_ACTIVE      ����   �$AP_AUTOMODE         �    �$AP_CHGAPONL         �   �$AP_COUPLED 1�������                                                                  �$AP_CUREQ 1������   T                                          	           	            	 ���                                          	           	            	 ���       �Handling      HT           	           	HTTHKY     	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ����$AP_CURTOOL      ����   �$AP_DO_CLEAN         �    �$AP_DO_CLENM  �������                                                                                                                          �$AP_DSPDRYRN         �    �$AP_HIDE  ������� @                                                                                                                                                                                                                                                                 �$AP_MAXAPP         �   �$AP_MAXAX          �    �$AP_PLUGGED      ����   �$AP_PRC_DSBM  �������                                  �$AP_PROC_DSB         �    �$AP_SEGF_CHK         �    �$AP_SEG_CHKM  �������                                                                                                                          �$AP_SELAP  ������� @                                                                                                                                                                                                                                                                �$AP_TOTALAX      ����    �$AP_USENUM  �������   �$ARG_STRING 1������� 
�MENUS             
MENU_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                I/O SIGNALS       Tryout Mode       Input Simulated   Output Simulated  OVERRIDE = 100    In cycle          Prog Aborted      Tryout Status     	Heartbeat         MH Fault          MH Alert            n                  n                  n                  n                  n                  n                  n                  n                  n                  n                TOOL              
TOOL_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                WORK              
WORK_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                POS               	POS_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                DEV               	DEV_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PALT              
PALT_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                GRIP              
GRIP_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                USER              
USER_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PREG              
PREG_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                �$ARG_WORD ?	�������  	$         	[         	]         	�          	�          �$ASBN_CONFIG �������           �$ASCII_SAVE            �    �$ATCELLSETUP 	�������%  OME_IO                               %MOV_HOME                              %MOV_REPR                                      �$AUTOBACKUP 
�������    FRA:\                                             '`                       �                 15/12/04 02:01:34         �                          �                          �                          �                            ��                                                                                                                                       ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      �  RA:\_BACKUP_\ATBCKCTL.TMP DATE.DT                                                                                                �$AUTOINIT         �    �$AUTOMESSAGE        �   �$AUTOMODE_DO         �   �$AUTOMODE_OV         �   �$AUTOPAUSPOS !��������  ( ?�?�ٿ2��Vv����U>2��7�SE@         )�                                    9�                                    I�                                    (O����������������������������(O����������������������������(O����������������������������(O�����������������������������$AUTOPPOSTSK  �������                              �$AUTOUPDTMOD         d�   �$AXIS_COUNT 1������   �  � 	 �L {��!�<��4HmȤ         	  1�| ~�; R�Z w�2 _Ȳ 6�� C�f         	                                      	  i�CN 0����o/p���vP�[         	                                 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXIS_METER 1������   �  P 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXSCRDCFG 1������  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �$BACKGROUND         �   �$BACKUP_NAME 	�������	BACKUP    �$BACK_EDIT 1������� 
 �%-BCKEDT-                              %FOLGE011                              �     ��%-BACKUP-                              �    �                        %-BCKEDT-                              ��%-BCKED2-                              %UP002                                      ��%-BACKU2-                                    �                        %-BCKED2-                              ��%-BCKED3-                              %                                       0��      %-BACKU3-                                    �                        %-BCKED3-                              ��%-BCKED4-                              %�                                      ���      %-BACKU4-                                    �                        %-BCKED4-                              ��%-BCKED5-                              %�                                      ���      %-BACKU5-                                    �                        %-BCKED5-                              ��%-BCKED6-                              %�                                      ���      %-BACKU6-                                    �                        %-BCKED6-                              ��%-BCKED7-                              %�                                      ���      %-BACKU7-                                    �                        %-BCKED7-                              ��%-BCKED8-                              %                                       ���      %-BACKU8-                                    �                        %-BCKED8-                              ��%-BCKED9-                              %                                       ���      %-BACKU9-                                    �                        %-BCKED9-                              ��%-BCKCRT-                              %�                                      ���      %-BACCRT-                                    �                        %-BCKCRT-                              ���$BCK_NO_DEL         �   �$BGE_UNUSEND         �   �$BLAL_OUT �������  �   �$BWD_ABORT         �    �$BWD_ITR_RTN         ��   �$BWD_NONSTOP         �   �$CE_OPTION         �   �$CE_RIA_ID         �   �$CFCFG �������                      �$CF_PARAMGP 1�������                                                                                                     C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  D  D  D  D  D    C�  C�  C�  C�  C�  C�  D	� D  D"� D/  D;� DH  DT� Da  Dm� Dz  D�@ D�� D�� D�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�  �$CHECKCONFIG         �    �$CHG_PRI 1�������         ��������������������������������������������������������������������������������������������������������������������$CHKPAUSPOS 1�������  ,    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    �������������������������������$COCFG �������              �$CO_MORGRP 2�������  �   IC4  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  �$CO_PARAMGRP 2�������  ,       ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�  �$CPCFG ������          a�-                                                                                   
                                            ����                @                                 �`        �$CPDBG ������        )cpmidbg                                      �   �  :�  -|  -}       )cpmpdbg                                      �     �  j  k       )midbg                                        �     �  �  �       )mpdbg                                        �     �             )mgdbg                                        �     �   N   O       )mfdbg                                     ���������                    )ud1:                                              �$CPDBGDEF ������       )ud1:cpdbgbuf.txt                             �                    �$CP_L64FIX ������                                                                                                                                                                                                                                                                                                                                                                                                                                               �$CP_MCRGRP 2������     d   d   d   d   d   d   d   d   d   d   d   d�$CP_MORGRP 2������  �                 @���CH  BH   	 B��B��\B�#rB�c�C�C-x�D         	 C���D!7�C�d}Dxz�D_`	D\�5FXT�         	 Fɛ�F�9�F��Fa��FF%�F[bJH/{?        ?�                              CH  BH   	                                      	                                      	                                     ?�                              CH  BH   	                                      	                                      	                                     ?�                              CH  BH   	                                      	                                      	                                     ?�         �$CP_PARAMGRP 2 ������ <                       |  �     �  x    	 C>  C*  C0  C�  Cp  D>  E�           	 D>  D��D{l�E�  D�  Em� Gj`          	 D�  Dl)E3� F�  E��fE��fH|         ?�  >�33 ;��?   ?�         n   @   @�   5�@   @   ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    �������$CP_RSMOFST ������                  �$CP_T1_MODE !������     G   
?@      ;��
                                               �$CP_TESTDEF ������           �$CRCFG "�������                             C4  A�             �   x   A�  Cz  B�  CH  B�  CH  C  @�     -       :d�
�$CRI_CFG #�������   �$CRT_DEFPROG %�������%�                                      �$CRT_INUSER         �    �$CRT_KEY_TBL  ������   	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������͓�����������������������������耇���������������������$CRT_LCKUSER         �    �$CRT_USESTAT         �    �$CR_AUTO_DO        ��    �$CR_INDT_ENB         �   �$CR_T1_DO        ��    �$CR_T2_DO        ��    �$CSTOP         �   �$CSXC_PARAM 2$������ 
 8
SONY XC-56                    �  �@���?�     ( АSONY XC-HR50                  �  �@���?�     ( АSONY XC-HR57                  �  �Aff?�     ( А�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �$CTRL_DELETE         �   �$CT_POPUP             �    �$CT_QUICKMEN         �    �$CT_SCREEN �������kcsc  �$CT_USERSCRN �������c_sc  �$CUSTOMMENU 1%������  <               %                                                          %                                       ���               %                                       ����              %�                                      ����              %�                                      ���Start SM Comm %IBSCMANS                              ���End SM Comm   %IBSCMANE                              ���User Cancel   %UCANCACT                              ���
User Reset    %URESACT                               ����              %�                                      ����              %�                                      ����              %�                                      ���Zange         %ZG_MENUE                              ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���VAG_KONFIG.   %VW_MENUE                              ����              %�                                      ���VAG-Dateien   %DATEIEN                               ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���
Macro Step tt %MSK_STAT                              ���Wait Monitor  %SHTPEST                               ����              %�                                      ����              %�                                      ���CYCLE POWER   %PWDCYCLE                              ���
POWER DOWN    %	PWD_MAINT                             ����$CUST_MANUAL         �   �$CZCDCFG &�������            	                                              ?|(��$DBCONDTRIG         �   �$DBLOVRD_ENB         �   �$DBNUMLIM        d�   
�$DBPXWORK 1'�������                                                                                                                          �$DBTB_CTRL (�������                ���$DB_AWAYTRIG      GCP �=��
�$DB_AWAY_ALM         �    �$DB_CONDTYP         �   �$DB_DBG 1)�������  , 
               	�   �   �  	|  	{   �     
                                        �$DB_MINDIST      GCP �@�  �$DB_MONTIME        ��  ��$DB_MONTYP         
�   �$DB_MOTNEND         �   �$DB_RECORD 1/�������  �                        G�O�G�O�   #            t/��t/�G    t/��  XECUTING

 ����                                                                  G�O�                                    G�O�G�O�   %            t/�Kt/�    t/�qEXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   &            t/��t/�w    t/��EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�               t/�"t/��    t/ިEXECUTING

 ����                                                                  G�O�                                    G�O�G�O�               t/�3t/��    t/��EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   S            t/|
t/}7    t/|iEXECUTING

 ����                                                                  G�O�                                    G�O�G�O�                                  XECUTING
  ����                                                                  G�O�                                    G�O�G�O�                                  XECUTING
 �����                                                                  G�O�                                    G�O�G�O�                                  TOPPING
                                                                       G�O�                                    G�O�G�O�                                  CANCELLED
                                                                       G�O�                                    G�O�G�O�                                                |[�                                                                G�O�                                    G�O�G�O�                                                p��                                                                G�O�                                    G�O�G�O�                                                                                                                   G�O�            �$DB_TOLERENC      B�  �=L���$DCSS_DEVICE 10������                                                                                                                                                                                                                            �$DCSS_LS 11������                                                                                                                                                                  �$DCSS_PARAM 2������                 �$DCSS_RBT 24������ 8 
 <                  Cπ       ¤  �H     �� �H                       Ck        ��  ��  �\  �g@ ��  �\                    C�        ��  B   �p                                B�                â�         ĸ`                   C1            �  ��      �             c                                                     c                                                     c                                                     c                                                     c                                              C��Dz  C��Dz   	 B��Aə�AU��A���A���B.��             	 B�  B�  B�  B�  B�  C>               	 B(  B��B��B[33BD��B�ff             	 B�  B�  B�  B�  B�  C>               	  �a� �G� X( X�� Q�� vy� j�x             
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                         �$DCS_CFG 5�������          dMC:\DCSL%04d.CSV                     c                   �    A   A   CH  Cz                                                                                �            �   �   �   �   �   �   �            �`iMU��    �$DCS_CRC_OUT 6�������                  �$DCS_C_FSI ?������ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_FSO ?������ P �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_RPI ?������  �                      �                      �                      �                      �$DCS_C_RPO ?������  �                      �                      �                      �                      �$DCS_SGN 7�������h��%12-JUN-24 17:02   ���04-DEZ-15 02:02            W"kJW"kJI$�H<6�                    h��%N��h�6%ZX�_                  �$DCS_VERSION �������V3.3.2            �$DEFLOGIC 18�������  	�          ���	�          ����	�          �����$DEFPROG_ENB         �   �$DEFPULSE         ��   �$DEF_ACCLIM        ��   ��$DEF_WRSTJNT         �����$DEMO_ENB            �    �$DEMO_INIT 9���������������� ���$DEMO_OPT_SL ?	������   � 
 	R575      	R745      	R746      	R747      	R750      	R751      	R752      	�          	�          	�          �$DEMO_OPT_TO  ������   � 
                                         �$DEV_INDEX         d�   �$DEV_PATH A�������A\KJLTVR411670R01\ 1670R01\ NGLISH\  EPASSAR TRAJETORIAS\          �$DHCP_CLNTID ?�������  �                  �                  �$DIAG_GRP 2>������ �    	 E�  F,D F,D E(p E(p D�               	 B�  B�  B�  B�  B�  B�               	 B�  B�  B�  B�  B�  B�               	 CeEC�� C�� CG�SCEZXB�Gm            f362 678901234567890          �  A���A�=qA�A�33A�z�A��A��RA���A�=qA���                  @�  A   Ap  A�  A�  A�  B  B   B4                        ������       
  A�A�{A�=qA�=qA�{A�A�G�Aď\A��A�Q����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A�=qAυAʣ�AŮA��\A�G�A��A�ffA���A��R���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A_�AZffAUG�AO�
AJ=qAD��A>�RA8��A2ffA,  ���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A`��A[�AV{AP��AK
=AE�A?33A8��A2�\A+�
���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A��
A��RA
=Axz�AqAj�RAc�A\Q�AT��AL�����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
 	 A�z�A�{A��\AJ=qAK
=Aq             	 =�G�=�G�=�G�>8Q�>8Q�>8Q�             	 8��b8��b8��b7�Ŭ7�Ŭ7�Ŭ             	 @ʏ\@ʏ\@ʏ\@�p�@�p�@�p�              @�  Ah  A�       	 <�C�<�t�=�P=�hs=�t�=��P             	 ;��
;��
;��
<#�
<#�
<#�
                 �?+ƨC�  <(�U     4 	 @���@���@���@���@���@���            A@     ?     	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	 ?Tz�?Tz�?Tz�?#�
?#�
?#�
             	 ��G���G���G���G���G���G�             	 B   B   B   B   B   B                	 Bx  Bx  Bx  A�  A�  A�               	 Ce
C�� C�� CG�{CEY�B�G�             	                                	   p  '  �  p  p  p             	 Ap  Ap  Ap  Ap  Ap  Ap               	 ED  E�� E�� D�� D�� DD               	                                         8��� 6b:��l��Y==�h?�6��?���hæ|,E�V�D�   �        	                                      	                                      	                                  æ|,E�V�D�B� !:�e�C3��     	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                 �$DICT_CONFIG ?�������          eg      ���$DISTBF_TTS         
�   �$DISTBF_VER        
�   �$DMAURST         �    �$DMSW_CFG @������               �$DOCVIEWER A������     	 ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  �$DPM_CFG B������                          
        �$DPM_SCH 2H������ 
�   Schedule 1            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 2            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 3            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 4            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 5            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 6            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 7            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 8            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 9            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 10           �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz  �$DPM_SIM 2I������                                                                                                                                                          �$DRC_CFG J�������!�                                  !�                                  !�                                  !�                                  !�                                     �$DSBL_FAULT K�������        �$DSBL_GPMSK         ��    �$DTDIAG L������            UD1: 678901234567890                         P                                                                                                                                                                                                                                                                                                                                              �               @   �$DTRECP L������            
UD1:                                          P                                                                                                                                                                                                                                                                                                                                              �               @   �$DUMP_OPTION  �������    �$DUTR_CFG      ����   �$DUTR_CPMES      ����   �$DUTY_TEMP  È�3B�  �A�  �$DUTY_UNIT         �    �$DYN_BRK M�������        �$ED_SIZE    '   �  x �$ED_STATE         �    �$EMGDI_STAT      ���     �$ENC_STAT 1N������  �                                                                     
                 d                                                                                                                                                                                                                                                                                                                                                                                                                                 ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        �$ENETMODE 1O�������                                            �$ERROR_PROG %�������%�                                      �$ERROR_TABLE  �������  �������������������������������������������������������������$ERRSEV_NUM       ��   �$ER_AUTO_ENB         �    �$ER_NOAUTO P�������          *�  *�  *�  *�  *�  +                                                        �$ER_NOHIS         �    �$ER_NO_ALM 1Q�������  �         *�  *�  *�  *�  +                                                                                                                                            �$ER_OUT_PUT 2R�������    @�                ����$ER_SEV_NOAU  �������                 �$ETCP_VER !�������!�                                  �$EXTLOG_REQ        ��    �$EXTLOG_SIZ        ��    �$EXTSTKSIZ        ��  ��$EXTTOL      Dz  �A   �$EXT_BWD_SEL         �    �$EXT_DI_BWD S�������                  �$EXT_DI_STEP S�������                  �$E_STOP_DO        ��    �$FACTORY_TUN         d�    �$FDR_GRP 1T������  d 	                             	 �[���.��FT&hB�( � ��� ��� 	                                      	     Bn�(B��@9LA��r@@�J             	     B]a�BuO�    A���                 	                                      	                                      	 A�A�5A��g@�H@��@��0             	 �|���hi�W���������/����             	 <��>    =(��<`�><��>                 
 GG�BuO�=(��    A��                         �                 	                                      	                                      	 C��NC��NC��NB�ƈB�ƈB�ƈ             	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	 E�� F@ F@ E�� E�� E��              	 OHcGPPL�uSL�uSK�y
             	 ?�  ?�  ?�  ?�  ?�  ?�               	 :G:�:G:�:G:�9{��9{��9{��             	 �2�y �������� 2��*Xou:         	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FEATURE U������   HandlingTool          ����English Dictionary    ����Multi Language (GRMN) ����4D Standard           ����Analog I/O            ����Angle Shift           ����Auto Software Update  ����Automatic Backup      ����Background Editing    ����Camera I/F            ����CnrRndImp             ����Common calib UIF      ����Condition Monitor     ����Control Reliable      ����Data Acquisition      ����Diagnostic log        ����Document Viewer       ����Dual Check Safety UIF ����Enhanced User Frame   ����Ext. DIO Config       ����Extended Error Log    ����Extended User Frames  ����External DI BWD       ����FCTN Menu Save        ����FTP Interface         ����Group Mask Exchange   ����HTTP Proxy Svr        ����High-Speed Skip       ����Host Communications   ����Hour Meter            ����I/O Interconnect 2    ����Incr Instruction      ����KAREL Cmd. Language   ����KAREL Run-Time Env    ����Kernel + Basic S/W    ����License Checker       ����LogBook(System)       ����MACROs, Skip/Offset   ����MH Core               ����MechStop Protection   ����Mirror Shift          ����Mixed logic           ����Mode Switch           ����Motion Diag. Core     ����Motion Optm. Core     ����Motion Profiler       ����Motion logger         ����Multi-Tasking         ����PCM function          ����Position Registers    ����Print Function        ����Prog Num Selection    ����Program Adjust        ����Program Shift         ����Program Status        ����Program Viewer        ����RDM Robot Discovery   ����Remote Conn Standard  ����Robot Servo Code      ����SNPX basic            ����Shift Library         ����Shift and Mirror Lib  ����Socket Messaging      ����TCP Auto Set          ����TCP/IP Interface      ����TMILIB Interface      ����TP Firmware           ����TP Menu Accounting    ����TPTX                  ����Telnet Interface      ����Tool Offset           ����Torque Simulator I/F  ����Touch Panel           ����Trouble Diag. & Prev. ����USB port on iPendant  ����Unexcepted motn Check ����User Frame            ����VCalibration Common   ����Vision Core           ����Vision Library        ����Vision SP CSUI        ����Vision SP CSXC        ����Web Plus              ����Web Server            ����Web Svr Enhancements  ����iPendant              ����iPendant Grid Display ����iPendant Setup        ����iRCalib. Standard     ����iRCalibration AAVM    ����Independent Axes      ����Independent Axes      ����Independent Axes      ����R-2000iB/185L         ����Ascii Program Loader  ����Ascii Upload          ����AutoMode TP operation ����Basic Remote TCP      ����CE Mark               ����CPRUT                 ����CRT/Keyboard Manager  ����Cntrl stop by E-Stop  ����Collision Guard       ����Collision Guard Pack  ����Constant Path         ����CornerDistance        ����Cycle Time Priority   ����DCS Joint Speed check ����DCS Safe I/O connect  ����DHCP                  ����Domain Name Serv.     ����Dyn Path Modifier     ����Enhanced Dry Run      ����Error Code Output     ����Ext Path Optimization ����Extended Axis Control ����External mode select  ����FRL Params            ����HMI Device (SNPX)     ����Integrated PMC        ����Internet Conn/Custo   ����Jnt Position output   ����KAREL                 ����Multi-Group Motion    ����Operation logbook     ����PC Interface          ����PROFINET I/O          ����PROFINET Safety       ����PROGRAM/JOG Override  ����Password Protection   ����PathSwitch            ����SNTP Client           ����TCP SPEED OUTPUT      ����User Function         ����User Socket Msg       ����VAG Package           ����VAG servogun setup    ����VAG setup 3           ����Weaving               ����iRCalibration VAxis   ����64MB DRAM             ����64MB FROM               �Arc Advisor            trsAux Servo Code        r
!Cell I/O              INT Common shell          ay SCommon shell core     AD pCommon softpanel      " #1Common style select   x_loCorner Region         rsv\Cycle time Opt.       ductDCS Pos./speed common AD pDisp 2nd analog port  
PCVEMAIL Enhancements    e4.pEmail Client          fx_mEnhanced Rob Serv Req \trsEnhanced T1 Mode      roduExt weave sch         LOADExtended Axis Speed   c
PFunc stup             otn.OPT TP Ins            
! nPC Send Macros        ionReal Simple Syn.(RSS) PRINRequires CP            PosRobot Library Setup   AD pRobot Service Request " #1SMB Client            \etnSSPC error text       nompSoft Limit            -fleSpace Check           H549TCP Speed Prediction  -fleTCPP Extention        AD pTrack Instruction     F" #Tracking Softpart     \fx_VAG Software          fxuiistdpnl               oducVAG V8.x Customizatio LOADVAG EMZ & EQ Tools    ENDIFREU late Updates     .comUpdate VAG PMC        ete"Ascii Upload when arg ����Profinet and CD Setti ����*.pc protection and u ����DryR.Skip PWF,VAGBCK  ����Activate CD Setting   ����VAG Menu to Page 1    ����Implement Feedb.Tig/T ����Fix upper limit of GO ����To fix skip problem   ����Files Updated         ����Activate CD-PS-Impr   ����Diff.a.DryS.PN:FW-CHK ����Diff.a.DryS.PN:FW-CHK ����CD:Fix SSTEP and BWD  ����Fix.Er.after 8xVag_C. ����Update several Issues ����Enh.Alloc.Mem.CD-Mot  ����To fix skip problem I ����Fix Err.Karel Var.Scr ����Fix DCS FB_CMP alarm  ����Fix overwr.VAG FUNC-M ����Restore Optimizations ����Fix.Karel User n.save ����ZIP cmd.er.handl.impr ����Restore Optimization  ����VAG Sign Off Function ����ATSHELL Heartbeat Opt ����No Outp.On/Off w.SRVO ����Fix-PS strt move away ����GunM.DO.Prot.Gen.Opt. ����Fix iPend.scrn freeze ����P381+Investig.Patch   ����Fix ABC Over Run      ����Over.disp.unexp.clear ����Inv.probl.about PGPX  ����Res.TCPspdoutVar E-St  k|Fix ABC Ov.load MSTP  pclsModification of iRCal ripcUnzip Inst+Improv.    roduFix PGPX OX-144 probl 
PCVEnh.DryRunP.Canc/Res  nopaFix OS144 Motn-UserCa hgriImprove VAG-Backup     proImprove VAG-Backup    c
P�                      mhse�                      \mhg�                      AD p�                      pc
�                      \mhv�                      t\mh�                      OAD �                      t.vr�                      !
!�                      l
!�                      Load�                      art �                      emov�                      LOAD�                      "FCT�                      emov�                      oduc�                      CVLO�                      orc.�                      val\�                      duct�                      LOAD�                      pc
�                      mr_w�                      remo�                       pro�                      
PC�                      t_to�                      emov�                      prod�                      
PCV�                      lwt.�                      val\�                      duct�                      D pr�                      
PC�                      _pre�                      d
!�                      ingu�                      
PR�                      ine �                      
TXP�                       "SI�                      siad�                      fd
�                      nse �                      G H5�                      SPLG�                       II)�                      plug�                      ealp�                      isp �                      ORDE�                      760 �                      Part�                      r760�                      AD p�                      
PCV�                      lt.p�                      sptk�                      \r76�                      .fd�                      le E�                      RINT�                      le E�                      �	��                      ct\j�                      rodu�                      AD p�                      PCVL�                      
PC�                      vr
�                      576.�                      j
!�                      INT �                       Hei�                      LOAD�                      OF" �                      \tho�                      t\j5�                      prod�                      VLOA�                      pc
�                      bwd.�                      ER R�                       RBW�                      
TXP�                       "RW�                      rbwd�                        ! �                       - R�                      ORDE�                      "Loa�                       Lib�                      oduc�                      VLOA�                      d1.p�                      !
!�                      
IF �                      Load�                      t II�                      e\aw�                      prod�                      1
P�                      dump�                      
! �                      d Eq�                      587 �                      E (R�                      II) �                      ld2\�                      duct�                      NDIF�                      63.f�                      ORDE�                      663 �                      "
P�                      w2tg�                      
! �                      
IF �                      ng J�                      ) "�                      cutx�                      722\�                      duct�                      AD p�                      
PCV�                      t1.p�                      wvcu�                      \j72�                      rodu�                      LOAD�                      c
P�                      vrcf�                      2\wv�                      ct\j�                       pro�                      CVLO�                      .pc�                      �[�                      TXPL�                       "FR�                      syrs�                      Tert�                      ENDI�                      amp.�                      RDER�                      INT �                      p, P�                      ct\s�                      XPLO�                      m "S�                      p.fd�                      mit�                      641 �                       H60�                      06 H�                      H629�                      7 H7�                      612 �                       H62�                      99 H�                      H663�                      MT (�                      TXPL�                      "FSL�                      lmt\�                      d
!�                       Uti�                       H89�                      Posi�                      I) "�                      os "�                      d
!�                       Axe�                      NT "�                       Axe�                      rodu�                      ENDI�                      ex.f�                      IF O�                      g H6�                      t II�                      ndex�                       ! a�                      Comp�                      ER C�                      adin�                      e, P�                      ct\c�                      a.fd�                      Envi�                      X H8�                      CFLX�                      rt I�                      lx\c�                       pro�                      CVLO�                      pc
�                      870.�                       ORD�                      H870�                       "
�                      r "R�                      d
!�                      ion �                       H82�                      997 �                      art �                      997\�                      D pr�                      F  !�                       M-1�                         �                      90" �                      \cle�                      rodu�                      
PC�                      m.pc�                      li_v�                      j590�                      uct\�                       pro�                      CVLO�                      .pc�                      02.p�                      e_no�                      0\wr�                      j590�                      ct\j�                      oduc�                      AD p�                      VLOA�                      
PC�                      ing.�                      \ext�                      j590�                      oduc�                      OAD �                      
PCV�                      rd.p�                      amdp�                      \j59�                      .fd�                      ppli�                       J59�                      Comm�                       "
�                      pc "�                      \cma�                      OAD �                      
PC�                      it.p�                      ! is�                      r
!�                      Load�                      , Pa�                      t\is�                      PCVL�                      .vr�                      
! i�                      r
!�                      Load�                      , Pa�                      t\is�                      CVLO�                      r
E�                      isds�                      g
!�                      Load�                      ing,�                      duct�                      
PC�                      s.vr�                      
! j�                      IF O�                      g J6�                       "
�                       "SV�                      41 H�                      OAD �                      S" #�                      fd
�                      h fo�                      2
P�                      oTor�                      
TX�                      r.pc  H552  oducH521  tsrsH532  CVLOR782  ct\jH550  pushJ614  LOADATUP  \j88J545  .pcJ616  ! j8VCAM  
! CRIM   - ECUIF  SnifJ628  IF OCNRE  9 R6R631  J598RSCH  88 JDOCV  NT "DCSU  R659J604  et SEIOC  PartR542  TXPLR696  uct\ESET  hcsnJ516  #1
J716  prodMASK  f\hcPRXY  NDIFJ627  f.fdHOCO  993.J513  alibJ542  MCalJ510  ORDEJ650  669J539  LoadH510   (iRLCHK  ion OPLG  art J503  XPLOMHCR  ct\jMCSP  mg "J506  
PCJ554  oducMDSW  cmg_MDCO  PCVLOPCO  uct\MPRO  g_exR637  VLOAJ600  t\j9PCMF  lib.J514  OAD J507  j993J515  .pcJ517   proJ505  3\vtPRST  
PCVJ697  ductFRDM  recpRMCN  LOADH930  \j99SNBA  r
ESHLB  j993SMLB  ! cvR636  VisiJ520  ommoHTCP   ORDTMIL  R669R789  90 JTPAC   R81TPTX   "LoTELN  VT (J509  CP cJ882  art R781  CVLOJ958  ct\cJ957  initUECK  LOADUFRM  \cvvVCCM  t.pcVCOR   ! cVIPL  !
!CSUI   - ACSXC  t (pWEBP  
IFHTTP  576R626  LoadCGTP   (ABIGUI   (pcIPGS  rt IIRCL  PLOAJ888  t\r5H895  i "AH895  
PCVH895  ductH613  ui.vR796    ! R507  
!
J698  d - R657   PxCJ618  !
IJ858  J896J535  "LoaJ570  6 (IR534  PxC J684  art R663  XPLOR748  ct\jJ523  ps "J555  
TXJ568  oducR526  tibsJ755   #1R739   proJ985  6\ibJ527  NDIFJ829  .fdJ518  dr.fJ569   MotR651  
!R553  R DMJ760  H798R558  99 HJ966   H87R632   "LoJ601  DR (J695  or DR641  rt IJ930  PLOAJ931  t\dmJ579  r "DJ541  
ENDJ693  dr.fR610  j932J694  sitiJ986  ordR648  RDERJ658  RINTJ653  g J9J656  tionJ504  d, PJ996  "
PD064  roduF064  pstrR666  
PCVSVMO  ductCLIO  tr_dR645  CVLOCMSC  ct\jCMSP  _dc2STYL  LOADR654  \j93CTOP  nd.pDCSC  AD pR528  932\JNN8  .pcJNN7   proORSR  2\psR680  c
PJ881  roduEXTS  pstrFCSP  
PCVOPIS  ductSEND  tr_sR679  CVLOCPRQ  ct\jRLCM  _wrtSRSR  LOADR677  \j93ETSS  py.pSLMT    ! J609  
!
J524  �*0TCPE  2\vtTOAW  
PCTRAK  oducFVAG  tmgrIPNL  CVLOVAG1  ct\jEZEQ  in.pUPD3  AD pPMC3  832\P137  c
PE001  roduE002  vtmuE003  CVLOE004  ct\jE005  s2.pE006  AD pP170  832\P171  c
PE007  roduRT22  vtprE008  PCVLE009  uct\P208  qpu2E010  LOADE011  \j83RT23  2.pcP213  D prP225  32\vP230  c
PP231  roduE013  vtvqP238  
PCVP244  ductE014  mofqP246  NDIFS300  .fdP275  58.fP276  T
!E015  ER JP381  NT "P477  J858P501   ParP525  
TXPP537  ductP333  zvsyE016  #1
P307  prodP576  \mnuP604  
PCVE018  ductP623  sy.vF001    ! F002  
!
�      d - �       Tor�      !
I�      R744�      "Loa�      4 (i�      Torc�      art �      CVLO�      ct\r�      elp.�      OAD �      r744�      .pc�       pro�      4\ir�      
PC�      oduc�      rtfl�      PCVL�      uct\�      kini�      VLOA�      t\r7�      in.p�      AD p�      744\�      pc
�      prod�      \irt�      c
E�      r744�      ! cv�      - iR�      for �      !
I�      VIRC�      00 J�       J91�      901 �      8 J9�      R730�      13 J�       R71�      738 �      INT �       VIR�      nect�      isn,�      ) "�       pro�      irc\�      .pc�      ! cv�      
!
�      d - �       Bin�      
!�      R J9�      T "L�      909 �      n Bi�      g, P�      "
T�      rodu�      bpfk�      #1
�       j90�      
! c�       - V�       VGF�       ORD�      J900�      12 J�       R68�      686 �      2 J9�      J840�      RINT�      g VG�      on S�      Part�      TXPL�      uct\�      pvgf�       #1�       pro�      gfs\�      .pc�       pro�      gfs\�      
END�      vgfs�      ! cv�      - Vi�      CCRG�      ORDE�      912 �      5 J9�      J904�      46
�      oadi�      (Vis�      CRG,�      ) "�       pro�      crg\�      CCRG�      VLOA�      t\cv�      rgtr�      VLOA�      t\cv�      rggt�      VLOA�      t\cv�      rgut�      VLOA�       ;�         �      1
P�      adin�      Remo�      or T�       II)�      OAD �      j941�      d.pc�       ! j�      !
!�       - V�      acki�      F OR�      
PR�      ding�      isua�      ng, �       "
�      prod�      \etv�      K" #�        ! �      
!
�      d - �      ogun�      !
I�      J653�      "Loa�      3 (V�      gun �      art �      CVLO�      ct\j�      ervo�      LOAD�      \j65�      1.pc�      D pr�      53\i�      pc
�      prod�      \vwe�      
IF�      656�      CVLO�      ct\j�      emz.�      F
I�      J656�      D pr�      53\v�      c
E�      DIF �      fd
�      4.fd�      etup�      F OR�      
PR�      ding�      AG s�      Part�      PCVL�      uct\�      ch_v�      VLOA�      t\j6�      _vw.�      F  !�      
!�      fd -�      up 2�      ORDE�      PRIN�      ng J�       set�      rt I�      VLOA�      t\j6�      _au.�      OAD �      j655�      u.pc�       ! j�      !
!�       - V�       3
�      DER �      INT �       J65�      etup�       II)�      OAD �      j656�      p.pc�      D pr�      56\p�      pc
�      prod�      \she�      
PC�      oduc�      ser_�      VLOA�      t\j6�      w.pc�      D pr�      56\v�      pc
�       J80�      
PCV�      duct�      io2b�      NDIF�      ER J�      LOAD�      \j65�      lt.p�      
EN�      656.�       fva�      AG S�      
!
�       FVA�      655 �      INT �       FVA�      oftw�      t II�      LOAD�      \fva�       "FE�      TXPL�      uct\�      ocm �      1
T�      rodu�      vwlo�      " #1�      D pr�      ag\v�      ENU"�      LOAD�      \fva�       "MO�      TXPL�      uct\�      skp �      1
T�      rodu�      vwne�      " #1�      D pr�      ag\v�      ARD"�      LOAD�      \fva�       "PF�      TXPL�      uct\�      lmn �      1
T�      rodu�      vwtt�      " #1�      D pr�      ag\v�      PPL"�      LOAD  H552      vwflH552        �H552         H552       (M-H552      t IIH552       proH552      c3 "H552      PLOAH552      74\pH552       #1H552      ductH552      c3.pH552      h774H552      hd.fH552      C
!H552      832H552      ing H552       iC,H552      
TXPH552      \nghH552      " #1H552      ghd.H552      r.fdH552      
!H552      33
H552      ng HH552      iC, H552      TXPLH552      ngdrH552       #1H552      dr.fH552      .fd H552      
!
H552      0
PH552      g H7H552      5, PH552      XPLOH552      710\H552      #1
H552      0.fdH552      fd -H552      
!
H552      1
PH552      g H7H552      0L, H552      TXPLH552      h711H552       #1H552      11.fH552      .fd H552      -30iH552      DER H552      "LoaH552      -500H552       ParH552      LOADH552      b\p5H552      
ENH552      fd
H552       - PH552      !
IH552      
PRH552       H68H552      5P, H552      TXPLH552      p70pH552       #1H552      0p.fH552      .fd H552      
!H552      84
H552      ng HH552      /15,H552      
TXPH552      \p70H552      " #1H552      70a.H552      s.fdH552      5S
H552      H686H552      dingH552      iA/1H552       "
H552      uct\H552      700"H552      ! p7H552      p70mH552      A/15H552      ER HH552      LoadH552      700iH552      II) H552      roduH552       "P7H552      F  !H552      
! pH552      00iAH552      ORDEH552      T "LH552      (P-7H552      rt IH552      D prH552      700 H552      NDIFH552      
!
H552      C-flH552      DER H552      "LoaH552      -fleH552      "
TH552      ct\hH552      AC" H552      prodH552      c "CH552      LOADH552      0\c5H552      
TXH552      t\h8H552      C" #H552      roduH552       "C3H552      OAD H552      \c4lH552      
TXPH552      \h82H552      " #1H552      oducH552      "CSLH552        ! H552      ! j6H552      r ReH552      �[H552      1
PH552      ct\jH552      
PCH552      t\j7H552      pc
H552      uct\H552      r.pcH552      oducH552      e.pcH552      oducH552      p.pcH552      oducH552      .pcH552      ductH552      fs.pH552      j726H552      83.fH552      n BiH552      
IFH552      
PRIH552      J783H552      Bin H552      t IIH552       proH552      actuH552      AD pH552      ikavH552      LOADH552      3\ikH552      CVLOH552      783\H552      
PCVH552      \j78H552      c
PH552      ct\jH552      .pcH552      ductH552      om.pH552      roduH552      nposH552       proH552      kindH552      AD pH552      ikli           LOAD           3\ik           CVLO           783\           
PCV           \j78           c
P           ct\j           .pc           duct           os.p           rodu           ckok            pro           prwo           AD p           ikpr           LOAD           3\ik           CVLO           783\           
PCV           \j78           c
P           ct\j           .pc           duct           ni.p           rodu           rial            pro           schn           AD p           iksl           LOAD           3\ik           CVLO           783\           
PCV           \j78           c
P           ct\j           .pc           duct           oc.p           j783           94.f           D OU�          ORDE�          T "L�          (TCP�          T, P�          XPLO�          694\�          " #1�          oduc�          p "T�          LOAD�          4\tc�            ! �          ! j5�          Spee�          
!�          24 H�          4 SL�          NT "�           (TC�          icti�           "
�          uct\�          "TCP�            ! �          ! rr�          Inte�          
IF �          PRIN�          RS1 �          ce V�          "
P�          ct\r�          c
P�          ct\r�          pc
�          1.fd�          �J��          ormm�          OAD �          \hi0�          VLOA�          39\n�          ENDI�          
!�           M-1�          IF O�          RINT�          27 (�          Part�          OAD �          \gnk�          
TXP�          \h82�          27" �          prod�          dgnk�           ! h�           h82�          /0.5�          ER H�          Load�          1iA/�          I) "�          oduc�          "M05�          AD p�          pfm0�          
PC�          t\h8�          pc
�          8.fd�          fd -�          
IF�          
PRI�          H813�          Part�          OAD �          \m11�          
TXP�          \h81�          13" �           h81�          741.�          S
!�          741�          ing �          3S, �          TXPL�          h741�           #1�          duct�           "GN�          OAD �          \pfm�          1
P�          ct\h�          c
P�          ct\h�          
EN�          fd
�           - M�          
IF �          PRIN�          742 �          Part�          OAD �          \m2s�          
TXP�          \h74�          CM" �          prod�          2sl �          CVLO�          742\�          CVLO�          742\�          DIF �          !
!�          -2iA�          RDER�           "Lo�          M-2i�          I) "�          oduc�          "M26�          AD p�          pfm2�          
EN�          fd
�           - M�          
IF �          PRIN�          744 �          Part�          OAD �          \m2h�          
TXP�          \h74�          44" �           h74�          701.�          A(B2�          RDER�           "Lo�          M-3i�          Part�          OAD �          \m36�          
TXP�          \h70�          CM" �          prod�          36a �          CVLO�          701\�          CVLO�          701\�          DIF �          !
!�          -3iA�          
IF�          
PRI�          H703�          203)�          
TX�           ��          PRIN�          629 �          P, P�          XPLO�          629\�          #1
�          uct\�          "H62�            ! �          ! h6�          0iA/�          ORDE�          T "L�          (M-9�          art �          AD p�          m92p�          TXPL�          h630�          P" #�          rodu�          2p "�          DIF �          !
!�          -900�          IF O�          RINT�          93 (�          , Pa�          PLOA�          93\m�          1
T�          ct\h�          H793�           ! h�           h79�          iB/7�          DER �          "Loa�          -900�           II)�          prod�          7 "M�          LOAD�          5\pf�          #1
�          5.fd�          fd -�          L
!�          796�          ing �          B/40�           "
�          uct\�          9B4"�           pro�          m9b4�          ENDI�          
!�           M-9�          
IF �          PRIN�          737 �          , Pa�          PLOA�          37\m�          1
T�          ct\h�          H737�           ! h�           h79�          0iA/�          ORDE�          T "L�          (M-2�          Part�          OAD �          \gzl�          
TXP�          \h79�          98" �           h79�          799.�          A/12�          DER �          "Loa�          -200�          rt I�          D pr�          dzl �          XPLO�          799\�          " #1�          799.�          9.fd�          175L�          R H6�          oadi�          000i�           II)�          prod�          7 "R�          LOAD�          9\pf�          #1
�          9.fd�          fd -�          0H
�          H610�          ding�          0iB/�          I) "�          oduc�          "R25�          AD p�          pfr2�          
EN�          fd
�           - R�          
!�          11
�          ng H  STD   B/15LANG   II)LANG  OAD STD   h611STD   21U"STD   LOADSTD   \h61STD    "H6STD     �STD   �[STD    - VSTD   ainiSTD   !
ISTD   CVSUSTD   12 JSTD    R68STD   686 STD   2 J9STD   J840STD   RINTSTD   g CVSTD   on TSTD   UIF,STD   ) "STD    proSTD   etu\STD   VISUSTD   PLOASTD   t\cvSTD   lmn STD   1
PSTD   roduSTD   u\vpSTD   c
PSTD   roduSTD   u\vlSTD   NDIFSTD   tu.fSTD   j512STD   ne TSTD   
!
STD    J51STD   945 STD   0
PSTD   adinSTD   LineSTD   g, PSTD   "
TSTD   roduSTD   lnlnSTD   " #1STD    ! jSTD   !
!STD   fd -STD   ostiSTD   F ORSTD    R81STD   021STD   LoadSTD    (iRSTD   ics,STD   ) "STD    proSTD   iag\STD   IRDGSTD   DIF STD   g.fdSTD   609.STD   ce CSTD   
IF STD   09 RSTD    R68STD    "LoSTD   09 (STD   eck,STD   ) "STD    proSTD   9\ssSTD   PC" STD   OAD STD   j609STD   
ENSTD   609.STD    etsSTD    SSPSTD   textSTD   ORDESTD   651 STD   1 R7STD   R683RBT   BI ARBT   NT "RBT   ETSSRBT   rrorOPTN  art OPTN  XPLOOPTN  ct\eOPTN  sspcOPTN  #1
OPTN   etsOPTN  !
!OPTN   - POPTN  aceOPTN  RDEROPTN  90 ROPTN   J94OPTN  945 OPTN  1 R7OPTN  J949OPTN  13 JOPTN  NT "OPTN  R641OPTN  erfaOPTN   II)OPTN  OAD OPTN  pcifOPTN  v.pcOPTN   ! pOPTN  !
!OPTN  .fd OPTN  l
!OPTN  ER IOPTN  
PROPTN  dingOPTN  stdpOPTN   II)OPTN  OAD OPTN  istdOPTN  vr.pOPTN  AD pOPTN  stdpOPTN  nl.pOPTN  AD pOPTN  stdpOPTN  st.pOPTN  DER OPTN  0 H5OPTN  OAD OPTN  istdOPTN  enk2DPND  IF
DPND   H52DPND  527 DPND  8 H5DPND  OAD DPND  istdDPND  ene2DPND  IF
DPND   istDPND  
!
DPND  fd -DPND  isorDPND  ORDEDPND  651DPND  LoadDPND   (ArDPND  r, PDPND  "
IDPND  ARCRDPND  74
DPND  prodDPND  v\awDPND  VS" DPND  F
IDPND  ARCRDPND  74
DPND  prodDPND  v\awDPND  VD" DPND  F
EDPND  awadDPND  
! oDPND  d - DPND  ns
DPND  DER DPND  1 R5CUST  
PRICUST  ing CUST  T TPCUST  rt ICUST  PLOACUST  �b�CUST   RRSCUST  551 CUST  1 R6CUST  J909CUST  30 JCUST   J94CUST  692 CUST  2 R7CUST  
PRICUST  ing CUST  b PlCUST   II)CUST  OAD CUST  webpCUST  ht "CUST  
PCCUST  oducCUST  s\hcCUST  NDIFCUST  lus.CUST   vcaCUST  amerCUST  
IFCUST  CAM CUST  0 H5CUST  H558CUST  CL CCUST   J87CUST  912 CUST  1 H5CUST  R685CUST  09 CCUST   R73CUST  913 CUST  C J8CUST  J888CUST  47
CUST  oadiCUST  (CamCUST   ParCUST  
TXPCUST  duct�      mncv�      #1
�      prod�      \etc�      S" #�        ! �      
!
�      d - �      alib�      
IF �      IF H�       H57�      558 �      L H5�      H574�      52
�      oadi�      (Com�      b UI�      II) �      AD p�      uif\�      CUIF�      DIF �      fd
�      iew.�      gram�      
!
�       J69�      590 �      6 H5�      H548�      74 H�      NT "�      J697�      m Vi�      rt I�      PLOA�      t\tp�      pvw �      1
E�      tpvi�      
! �      .fd �       Dia�      
!
�       MDC�      590 �      6 H5�      R765�      48 H�       R71�      021 �      INT �       MDC�      n Di�      , Pa�      
TX�      oduc�      nd\d�      GPT"�      IF  �      nd.f�      skmg�      cket�      ng
�      DER �      1 R5�      R651�      73 H�       J94�      549 �      O R7�      R641�      83 R�       RRS�      551 �      8 J8�      R710�      11 S�       R83�      949 �      3 J9�      
PRI�      ing �      cket�      ng, �       "
�      prod�      \tph�      M" #�        ! �      
!
�      d - �      Diag�      .
!�      ER J�       H59�      596 �      9 MD�      R818�      51 H�       S01�      552�      Load�       (Tr�      ag. �       Par�      
TXP�      duct�      dtrc�      #1
�      prod�      \sfm�      R" #�        
��         �         u�      T�EM�      ���$�       ��      �����      OST��      ?��      H573�      58 H�       H55�      583 �      9
P�       x�         �      716\�      HCHS�      PLOA�      t\j7�      p "P�      
PCV�      duct�      hs.v�      AD p�      716\�      
END�      16.f�      tcpi�      CP/I�      ace�      RDER�      41 R�       R65�      573 �      8 J9�      H549�      LN H�       SNB�      RCL �      C WE�      MDCO�      CO R�       R66�      818 �      3 R8�      R626�      55 R�       R61�      945 �      4 R5�      R540�      04 R�       RRS�      912 �      8 H5�      R648�      85 R�       R68�      902 �      6 J8�      R659�      92 R�       R58�      597 �      8 S0�      H552�      59 J�       R78�      689 �      9 PT�      J989�      47
�      oadi�      (TCP�      rfac�      II) �      AD p�      cpip�      "HCT�      XPLO�      ct\t�      cpp �      1
T�      rodu�      \tph�      G" #�      AD p�      cpip�      
PC�      oduc�      hcpg�      E
I�      R650�      ry
�       H52�       Sec�      PRIN�      tion�      ding�      CP/I�      ace,�      ) "�       pro�      ip\t�      CTC"�      LOAD�      \tcp�      p "H�      
TXP�      duct�      phcp�       #1�       pro�      ip\h�      PCVL�      uct\�      pg.v�        ! �      y
E�      Prim�      IF  �      fd
�      tcom�      ost �      atio�      F OR�       H54�      593 �      0 H5�      H558�      26 H�       HTC�      TTP �        ��      _T �       $M�      $VER�      EC �      1 R7�      R641�      12 R�       PRX�      526 �      0 R6�      JNN6�      38 R�       R53�      713 �      1 R7�      RRS2�      51 H�       J90�      688 �      6 R7�      J913�      40 J�        
��      �^��       !  �       �  �          �      ����      }��          �          �         H�          �      ����        
��      :PRO�      0\PR99    >_��$FEAT_DEMO U������   �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                            �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �            �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �                �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �$FEAT_DEMOIN         ��   �$FEAT_INDEX         ��   ��$FILECOMP V�������        �$FILESETUP2 W�������  �  N   N �$FILE_AP2BCK 1X������  �)MAKRO900.TP                               %MAKRO900                                 %MAKRO900                                  )MAKRO910.TP                               %MAKRO910                                 %MAKRO910                                  )MAKRO920.TP                               %MAKRO920                                 %MAKRO920                                  )MAKRO930.TP                               %MAKRO930                                 %MAKRO930                                  )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_APPBCK 1X������ 2 �)*.VR                                      %*                                         %                                           )*.PC                                      %FR6:*.PC                                 %                                           )*.TX                                      %FR6:*.TX                                 %                                           )*.FVR                                     %	FR6:*.FVR                                %                                           )*.STM .STM                                %FR:*.STM .STM                            %iPendant Panel                            )*.HTM                                     %FR:*.HTM                                 %                                           )*.GIF                                     %FR:*.GIF                                 %                                           )*.JPG                                     %FR:*.JPG                                 %                                           )*.JS                                      %FR:*.JS                                  %
JavaScript                                )*.CSS                                     %FR:*.CSS                                 %Cascading Style Sheets                    )
ARGNAME.DT                                %FR:\ARGNAME.DT                           %ARGNAME                                   )	PANEL1.DT                                 %FR:PANEL1.DT                             %iPendant Panel                            )	PANEL2.DT                                 %FR:PANEL2.DT                             %iPendant Panel                            )	PANEL3.DT                                 %FR:PANEL3.DT                             %iPendant Panel                            )	PANEL4.DT                                 %FR:PANEL4.DT                             %iPendant Panel                            )SHELL.VR                                  %SHELL                                     %�                                          )ZG_MENUE.VR                               %ZG_MENUE                                  %�                                          )
EINGABE.VR                                %EINGABE                                   %�                                          )SUMM_VAG.DG                               %FR:SUMM_VAG.DG                           %�                                          )TPE_STAT.VR                               %TPE_STAT                                  %�                                          )
TPEINS.XML                                %FR:\TPEINS.XML                           %Custom Toolbar                            )PASSWORD.DT                               %FRS:\PASSWORD.DT                         %Password Config                           )VAGCONF1.XML                              %FR:\VAGCONF1.XML                         %�                                          )EXTSERVO.VR                               %EXTSERVO                                  %�                                          )	IO_SET.DT                                 %FR:\IO_SET.DT                            %�                                          )VWEMZROU.VR                               %VWEMZROU                                  %�                                          )VAGBCKUP.VR                               %VAGBCKUP                                  %�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_DGBCK 1X������ ( �)
SUMMARY.DG                                %MD:SUMMARY.DG                            %Diag Summary                              )
CONSLOG.DG                                %MD:CONSLOG.DG                            %Console log                               )	TPACCN.DG                                 %	TPACCN.DG                                %TP Accounting                             )FR6:IPKDMP.ZIP                            %
IPKDMP.ZIP                               %TP Exception                              )MD:MEMCHECK.DG                            %MD:SUMMARY.DG                            %Memory Data                            �)MD:SHADOW.DG                              %MD:SUMMARY.DG                            %Shadow Changes                        �_�)	FTPLOG.DG                                 %MD:SUMMARY.DG                           %Comment TBD                           \+�)ETHERNET.DG                               %MD:ETHERNET.DG                           %Ethernet Configuration                    )MD:DCSVRFY.DG                             %MD:SUMMARY.DG                           %DCS verify all                        �s�)MD:DCSDIFF.DG                             %MD:SUMMARY.DG                           %DCS verify diff                       �s�)MD:DCSCHGD1.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �G�)MD:DCSCHGD2.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �G�)MD:DCSCHGD3.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �G�)UPDATES.DAT                               %FRS:\UPDATES.DAT                         %Updates List                              )
PSRBWLD.CM                                %FRS:\PSRBWLD.CM                          %PS_ROBOWELD                               )MD:SMTPLOG.DG                             %MD:SUMMARY.DG                            %SMTP/Email diag                       �&|)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_FRSPRT  �������    �$FILE_MDONLY 1X������    
 �)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_VISBCK 1X������ 
 �)*.VD                                      %FR:\VISION\DATA\*.VD                     %Vision VD file                            )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FMR2_GRP 1Y������� �C4  B�   	                             	 E�� F@ F@ E�� E�� E��              	 OHcGPPL�uSL�uSK�y
             	 ?�  ?�  ?�  ?�  ?�  ?�               	 :G:�:G:�:G:�9{��9{��9{��             	 A�  A�  A�  A�  A�  A�  A�  A�  A�  BH   	 C��NC��NC��NB�ƈB�ƈB�ƈ                	                                      	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	 =���=�L�<���=�(H>C�s>�I             	 :���:��;%�9޹p9��:���             	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FMR_CFG Z������� T                                                                                    �$FNO �������F174584             @�$FRM_CHKTYP  ����   ������$FROMCHK_MIN        ���  X�$FSSB_CFG [������                                                                           �$FTP_DEF_OW         �    �$FTP_DIRCOMP         �    �$FUNC_SETUP  �������                                                                                  �$GENOVRD_DO        �   �    �$GENOVRD_THR         d   �   d�$GENOV_ENB         �   �$GRAVC_GRP 1\������  �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            ��$GROUP 1b�������                       8�?�              ?�              ?�                  8���  ���.    ����3;�.?�  ���.?�  �;�.D=  Cr        C�  C>                                                             B�Q�               B�                                                                 8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   81�?�              ?�              ?�                  81�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  C�  C�                                                              �                  B�                                             �$GRSMT_GRP 1c�������      C�      C�      C�      C�  �$HOSTC_CFG 1d������ ��                  	FTP       �            �                          172.26.32.230                e                                                                                                       e�                                                                                                      172.26.32.230         e	cfg_fanuc                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �$HOSTENT 1e�������  P!�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !QUICC0                                  !172.26.32.90                      !QUICC1                                  !�                                  !QUICC2                                  !�                                  !ROUTER                                  !172.26.32.1                       !PCJOG                                   !192.168.0.100                     !CAMPRT                                  !192.168.1.10                      !CAMRTR                                  !192.168.1.10                      �$HOSTNAME !�������!KJLTVR411670R01RS--KU1            �$HOSTS_CFG 1d������ �Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                                     	SM                     �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                            �    �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �$HOST_ERR f�������                    �$HOST_PDUSIZ     ^  ��  >�$HOST_PWRD ?������   �  backup        guest         guest         guest         guest         guest         guest         guest         �$HSCDMNGRP 2g������� �      Z               K       	P01.03 8   	   6  �  �  A  �  .  "         	 �������W���x������`�������a         	   �  
b    �  �  8             	 ���6�����������x�������             	   N    	�  /    u             	 �����������M�����������             	   �  �  �  �  �  �               Z 	   6  �  �  A  �  .             	 �������W���x������`����                  d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                     �$HSCD_GROUP 2h������      	HSCD01.01         �                  �                  �              �$HSCD_QUPD         �   �$HSCD_UPDTYP  �������   �$HTTP_AUTH 1i�������  <!iPendant                          �                    !KAREL:*                           �                    !KCL:*                             �                    !VISION SETUP                      �                    !�                                  �                    !�                                  �                    !�                                  �                    !�                                  �                    �$HTTP_CTRL j�������                 
 %�FFF9E3                       FRS:DEFAULT               FANUC Web Server             
�$HTTP_PWRD ?������   �  �              �              �              �              �              �              �              �              �$HWR_CONFIG k�������  f                    �$IBGN_CFG l�������       2   @   <#�
<#�
<#�
BH  <#�
<#�
<#�
CH            4   <#�
        �$IBGN_DEV       ���   �$IBGN_ERRIO m�������                �$IBGN_EXDAT n������   �            �$IBGN_EXFLG            �    �$IBGN_FIL o�������                    �$IBGN_FTP p�������                    �  �	MERCATOR  	RECORD    	R_ACHS    	R_ISTW    IBGN  IBG   	SENSPS    TXT   999   	Keine 0                                     %IBSCRECS                               8�%IBSCRECE                               ��           �$IBGN_LMTN  �������                                                                                                                          �$IBGN_SBADR      ���   ��^�x�$IDL_CPU_PCT      B�   B�ȳ�$IDL_MIN_PCT      B�   =f��$IGNR_IOERR        ���   �$INPT_SIM_DO        ��    �$INTPMODNTOL         ��    �$INTP_PRTY        ��    �$IOLNK 1q�������                                                                                                                                  �$IOMASTER         �    �$IOSLAVE r�������    �$IO_AUTO_CFG         �    �$IO_AUTO_UOP         �    �$IO_CYCLE         �    �$IO_DEF_ASG 1s�������              d                     d                �   c                �   c                  
   c                  
   c                                                                                                                                                                                                                                                                                                                                                                                                                 �$IO_DEF_NUM     ����   �$IO_IPCHE         �   �$IO_RTRY_CNT      ����    �$IO_SCRN_UPD        ��    �$IO_UOP_CFG t�������    �������������������������$ISDT_ISOLC  �������                  �$J23_DSP_ENB  �����������$JOBPROC_ENB         �    �$JOG_GROUP 1u������� 8   d8�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8!�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d81�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8A�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                �$JOG_IN_AUTO      ����    �$JPOSREC_ENB         �    �$KANJI_MASK        ���    �$KAREL_CFG v�������          �$KAREL_ENB         �   �$KCL_LIN_NUM         �   �$KEYLOGGING  ����   d�   �$LANGUAGE �������ENGLISH       �$LGCFG w�������         ��   x  �  �  H  �   '0           �                     MC:\RSCH\00\                 �$LN_DISP x�������                                                    �$LOCTOL      Dz  �A   �$LOGBOOK y�������   d               d  X                                                                                                                                              	LOGBOOK            ��                                                �$LOG_BUFF 1z�������                    d                         d                                                                                                                                                                                                                                                                                                                                                                                   �$LOG_DCS |�������    =���                                        �������������������������������������������������������������$LOG_DIO 1}�������  ������������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ����������������������$LOG_ER_ITM  ������� d                                                                                                                                                                                                                                                                                                                                                                                                                 �$LOG_ER_SEV  �������   �$LOG_ER_TYP  �������                                                                                  �$LOG_REC_RST         �   �$LOG_SCRN_FL 1~�������    �                                                                                                                                                           �$LOG_TPKEY  �������                 �$LONGNAM_ENB         �   �$LUPS_DIGIT         �   �$LU_LOADPROG %�������%UP027                                 �$MAXUALRMNUM       ��   
�$MAX_DIG_PRT        �   �$MCSP ������                               d                �$MCSP_GRP 2�������  �   2     	     �  �                         	                                      	                                             	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                     �$MD_LDXDISAB  �����������$MEMO_APNAME ?������� 
 �              �              �              �              �              �              �              �              �              �              �$MISC 1��������  � 	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                         �$MISC_MSTR ��������    �$MISC_SCD 1�������� 
 � 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$MKCFG ��������                       �$MLTARM_CFG �������          �����������������������������$MLT_GRP_DO ��������         ��L��                                                                                                                                        �$MMETPU       ���    �$MNDSP_CMNT         �    �$MNDSP_MST ��������                                              �$MNDSP_POSCF         �   �$MNDSP_PRPMT         �   �$MNDSP_PSTOL 1��������  4@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�$MNSING_CHK         �    �$MODAQ_CFG ��������                             �$MODAQ_DEV 	�������	MC:       �$MODAQ_HSIZE  �������   ��$MODAQ_TASK %�������%$123456789 123456789 123456789 123456  �$MODAQ_TRIG 1��������  l������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ����������$MODAQ_TYPE      ����   �$MODEM_INF 1������� `)AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          �$MONITOR_MSG ?	�������   	EXEC1     	EXEC2     	EXEC3     	EXEC4     	EXEC5     	EXEC6     	EXEC7     	EXEC8     	EXEC9     	EXEC10    	EXEC11    	EXEC12    	EXEC13    	EXEC14    	EXEC15    	EXEC16    	EXEC17    	EXEC18    	EXEC19    	EXEC20    	EXEC21    	EXEC22    	EXEC23    	EXEC24    	EXEC25    	EXEC26    	EXEC27    	EXEC28    	EXEC29    	EXEC30    	EXEC31    	EXEC32    �$MOR_GRP_SV 1�������  ( 	 ?�ٿ2��Vv����U>2��7�SE@          	                                      	                                      	                                     �$MOTASK_DATA  �������    �$MPL_NAME !�������!Default Personality (from FD)     �$MRR2_GRP 1����  	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                                
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                   E@ E�` E�           	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$MRR_GRP 1�������  `     � �     � @D�  D�  ?�  ?�   �?   ?�      @T;gD�  D�                             ;�	l?�   	 ����X�    	 �X^ �,X� � � 	 K��K�CK�zK~o�K{GK�MF�N�         	                      	   �  �  �  �  �  �  �  �  � 	 ?�;g?��N?Ę	@
�@
�@T;gD�                   	 �Iۿ�
��������X����/           	 �4  �p  ���ô  ��  ô               	     ��Pտ�n    ��                 	                     �   �   � 	                                	   �  �  �      �    �  � 	                                      	  	'� �  �  I� �  �� #��         	 :�È:�È:�È:�È:�È:�È=���=���=��� 	  @ @ @ @ @ @  ��         	   �  �  �  �  �  �  L�          �    	                               	   ��  ��  ��  ��  ��  ��  N   ��  �� 	 @I�?��@{S�@��@�X@��E��          	 C4  B�  Ca  C�  B�  C�                  ��C9   	  � ���        	        } } H       	 B�  B�  B�  B   B   B   C             @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  I� �  �� #��         �   � :=              �   ?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  ?      �?            	  (   (   (   P   P   P            	             �?333       	 ;��;QaT;\��;��;�	�<$DA�D         	                       A0              ?�   �    ?fff  ?fff?@  ?&ff?    	 A�A�A�@�,@�,@�,            C9    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	     E�  E;�     E@ E�`              	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ��H�'#Gxo�F��=̳sƌ� A�           	                                                                                       A�  �?��                    ��  BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                      	                                    	     ?��                             	                                      	             ��@     �k               	 C�  D�` Ca                           	 ?��    ���?�ؿ��@I�             	 D/�CG33Ck�B�1B-v�=���             	 ÙE�ីW
�u                     	 ²B���  AX��Blz��X��                 	 ³
=Õ��ö�=BU(���  ��              	 K��JD��LUW�H�� I%K�AP               	 LUL =�L]��HP� H�R�AP               	 LTF�L%�J�
`H㞀H���A�               	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	     G�>                              	     C�ٚ                             	     Ć�                             	     CV��                             	                                      	 �                                   	                                      	                                      	 ( 	 �`��                    ��������� 	     �$rc                ��������� 	         3-NQ            ��������� 	             3��v        ��������� 	             ��v3�g�    ��������� 	             �!�;�%D93ҵ���������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	       )                             	                                      	                �                     	               8  t                 	                                      	                                      	                                      	 ( 	                             	                             	      9                      	                             	            O�                	            �e 3�             	                             	                             	                                 2 E@         E�`         E�          B��A   A�  C�  D  A   @�                                      �                                   Gr0 F� G�� D	� C�              �                                        E@         E�`         E�                                                                                      ?�  ?�              	                               
                                                                                                                                                                                                                                                                                          	     ��            �uD�Y      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$MSKCFMAP  �������                               �$MSKCONREL         �   �$MSKEXCFENB         
�    �$MSKEXCFFNC         
�   �$MSKJOGOVLIM         d�   d�$MSKKEY         �   �$MSKKEY_PANL             �$MSKRUNOVLIM         �   �$MSKSFSPDTYP         
�    �$MSKSIGN         �   �$MSKT1MOTLIM         d�   �$MSK_CE_GRP 1��������  \     	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                        �$MSQZ_EDIT      ����    �$MTCOM_CFG 1��������         
       
       
       
       
       
       
       
�$MT_ARC_ENB         �   �$MUAP_CPLENB         �    �$NOCHECK ?�������  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �$NO_WAIT_LN        ���   �$NUM_RSPACE  �������     
   
   
   
   
   
   
   
�$ODRDSP_ENB         �    �$OFFSET_CART         �    �$OFFSET_DIS         �    �$OPEN_FILES     
   ��   
�$OPTION_IO         �   �$OPTM_PRG %�������%$************************************  �$OPWORK ��������     �� �� ��       ���                         	 �                      �      ��$ORG_DSBL  �������                                  �$ORIENTTOL      C�  �A   �$OUT_SIM_DO        �    �$OVRDSLCT ��������    ������   
   
   
   
    �$OVRD_PEXE         �    �$OVRD_RATE         d�   �$OVRD_SETUP ��������     
 ����������������������������������������     
 �����������������������������������������$PARAM2_GRP 1���� 	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                                
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$PARAM_GROUP 1�gX�� `     � �     � @D�  D�  ?�  ?�   �?   ?�      C>  D�  D�                             ;�	l?�   	 ����X�    	 �X^ �,X� � � 	 H��Hޓ�H�33H��H�WH-��F�N�         	                      	   �  �  �  �  �  �  �  �  � 	 B�  B�  B�  B�  B�  C>  D�                   	 �4  �p  ���ô  ��  ô  �/           	 �4  �p  ���ô  ��  ô               	     �����lu�    ���                 	                     �   �   � 	                                	   �  �  �      �    �  � 	                                      	  	'� �  �  I� �  �� #��         	 =���=���=���=���=���=���=���=���=��� 	  @ @ @ @ @ @  ��         	   �  �  �  �  �  �  L�          �    	                               	   ��  ��  ��  ��  ��  ��  N   ��  �� 	 C4  B�  Ca  C�  B�  C�  E��          	 C4  B�  Ca  C�  B�  C�                  ��C9   	       ��        	        } } H       	 B�  B�  B�  B   B   B   C             @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  I� �  �� #��         �   � :=             �   ?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  ?      �?            	  (   (   (   P   P   P            	             �?333       	 ;��;QaT;\��;��;�	�<$DA�D         	                       A0              ?�   �    ?fff  ?fff?@  ?&ff?    	 A�A�A�@�,@�,@�,            C9    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	     E�  E;�     E@ E�`              	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                       A�  �?��                    ��  BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                      	                                    	     ?��                             	                                      	             ��@     �k               	 C�  D�` Ca                           	 ?��    ���?�ؿ��@I�             	 D/�CG33Ck�B�1B-v�=���             	 ÙE�ីW
�u                     	 ²B���  AX��Blz��X��                 	 ³
=Õ��ö�=BU(���  ��              	 K��JD��LUW�H�� I%K�AP               	 LUL =�L]��HP� H�R�AP               	 LTF�L%�J�
`H㞀H���A�               	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	     G�>                              	     C�ٚ                             	     Ć�                             	     CV��                             	                                      	 �                                   	                                      	                                      	 ( 	 �`��                    ��������� 	     �$rc                ��������� 	         3-NQ            ��������� 	             3��v        ��������� 	             ��v3�g�    ��������� 	             �!�;�%D93ҵ���������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	       )                             	                                      	                �                     	               8  t                 	                                      	                                      	                                      	 ( 	                             	                             	      9                      	                             	            O�                	            �e 3�             	                             	                             	                                 2 E@         E�`         E�          B��A   A�  C�  D  A   @�                                                                          Gr0 F� G�� D	� C�                                                                                                                                                                       ?�  ?�              	                               
                                                                                                                                                                                                                                                                                          	     ��            �uD�Y      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$PARAM_MENU ?�������  DEFPULSE              	WAITTMOUT             RCVTMOUT              SHELL_WRK.$CUR_STYLE  SHELL_WRK.$CUR_OPTA   SHELL_WRK.$CUR_OPTB   SHELL_WRK.$CUR_OPTC   SHELL_WRK.$CUR_DECSN  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PASSREL_ID      ���   �    �$PAUSE_PROG %�������%�                                      �$PCCRT         �    �$PCCRT_HOST !�������!PCCRT                             �$PCTP         �    �$PCTP_HOST !�������!PCTP                              �$PC_TIMEOUT      ����   �$PGDEBUG  �������    �$PGINP_FLMSK      ����    �$PGINP_FLTR      ����   �$PGINP_PGATR  �������                     �$PGINP_PGCHK      ����   �$PGINP_TYPE ?������  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PGINP_WORD ?	�������  	FOLGE     	UP        	MAKRO     	SUCHL     	MAKROSP   �$PGTRACECTL 1�������� 
   � �   � �                                         �$PGTRACEDT Q�������� 
D � 	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  	� c  	� d  	� e  	� f  b   ��    J   J   J   b   b   b   	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  	� c  	� d  	� e  	� f  b   ��    �   ��    	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4   � 
 �  
 �  
 �  
 �  
  	S   

   

   

   

   

   

   

   

   

 	  

 
  

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

   

    	S   	S   	S 	  	S 
  	S   E   E   E   E   E    E !  E "  
�   
�   
�   
�   
�   
�   E $  
�   
�   
�   
   
   
   
   
   
   
   
   
 	  
 
  
   
   
   
   
�   
�   
�   
�   E &  
�   
�   
�   
�   
�   
�   ��    J   J   J   b   b   b   	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  	� c  	� d  	� e  	� f  b   
 �  
 �  
 �  
 �  
 �   � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    �$PGTRACELEN       ��   ��$PGTRACE_UP ��������   ����$PG_CFG ��������       ����                                                     �$PG_DEFSPD ��������  �     ��$PING_CTRL ��������      8       �$PIPE_CONFIG �����������                   �$PLID_CFG ��������   �$PLID_GRP 1������� �   C8���V    A�
=G� G�L�F�( A�  D	�          �   d      d      d   d   d   d         � 	                                    	                 ´  ´               	                 B�  B�               	                 ´  ´               	                 B�  B�               	                 B�wB<h�             	                                      	                 <,1<,1             	                                      	                                      	                                      	                 <,1<,1             	                                      	                                      	                 Dz  Dz                      
 C
��A�;����>AU)�E��3H���H�|�                     	                                      	                                      	                                      	                                      	                 >V�0>Wj             	                                      	                                      	                                        !    
V7.10beta1         @�@_\)@0��C9    C�C�B���  D�  D�  D0�   D�  D�� Df� C9  A�  B�  C9  C>  Ap     B�  B�  B���C;��BffB33Be33B$  B$  B$  B��BffB4��ºC�º݋��     ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ����$PLID_KNOW_M         �   �$PLID_SV ���������        
                                                                                  	                                      	                                        d      d   d    �$PLIM_GRP 1��������  lC9   	       ��        	        } } H       �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���$PLMR_GRP 1��������  T        B�  B�  C9      Cf   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�              �$PLST_GRP1 1�������� 
 0Vacia             B�Q�A'�YyA*�)    H\H��hLlena eza         C
��A�;����>AU)�E��3H���H�|��                  C9                          �                  C9                          �                  C9                          �                  C9                          �                  C9                          �                  C9                          �                  C9                          �                  C9                          �$PLST_GRP2 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP3 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP4 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP5 1��������  0�                  �<                         �$PLST_GRP6 1��������  0�                  �<                         �$PLST_GRP7 1��������  0�                  �<                         �$PLST_GRP8 1��������  0�                  �<                         �$PLST_GRPMAD        �   �$PLST_PARNUM  �������                              �$PLST_SCHMAD         �   
�$PLST_SCHNUM         �   
�$PLST_UPDNUM  �������                          �$PLS_CMP_LIM  ����  '�   �$PLS_ER_CHK  ���� ���    �$PLS_ER_LIM  ����  '�   �$PLS_ER_RST         �    �$PL_MOD         �   �$PL_MOD_ST         �   �$PL_RES_G1 1�������� 
  B�Q�C��C��C�/}I}�I}�H�5�   C
��DF�DF�C���I)V�I)V�If�                                                                                                                                                                                                                                                           �$PL_RES_G2 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G3 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G4 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G5 1��������                                  �$PL_RES_G6 1��������                                  �$PL_RES_G7 1��������                                  �$PL_RES_G8 1��������                                  �$PL_RES_V 1�������   �  �^�`�^��]���]���$PL_THR_INRT         d�   d�$PL_THR_MASS         d�   Z�$PL_THR_MMNT         d�   Z�$PMON_QUEUE ��������       �      �$PM_GRP 2�������  4      A�  @�                    B�           �$PNS_CUR_LIN        ���    �$PNS_END_CUR         �    �$PNS_END_EXE         �    �$PNS_NUMBER        ���    �$PNS_OPTION         �   �$PNS_PROGRAM %�������%PNS                                   �$PNS_TASK_ID        ���    �$POCFG ��������                                      �$PODATA_GRP 1�������� @  r>   . 2 �����*�����*�����*�����*����	I	I	I	I	I	I	I	I	I	I	I	I	I	I	I	I	I	I���* 2       
      
      
      
     O O O O O O O O O O O O O O O F O O    
 2                                                     �>    2 ���	I	I	I	I	I	I	I	I	I	I	I	I	I
�	I	I	I	I	I00	I	I	I	I������*������*�����**� 2     O O O O $ O O O   O O O  O O O O O  	 C D O O           3          	  2                                                     �>    2 ���	I	I	I	I	I	I	I	I	I	I	I	I	I
�	I	I	I	I	I00	I	I	I	I������*������*�����**� 2     O O O O $ O O O   O O O  O O O O O  	 C D O O           3          	  2                                                     �>    2 ���	I	I	I	I	I	I	I	I	I	I	I	I	I
�	I	I	I	I	I00	I	I	I	I������*������*�����**� 2     O O O O $ O O O   O O O  O O O O O  	 C D O O           3          	  2                                                   �$POINFO_GRP 1�������� �     �                                                                                                                                                                                                                                                                                                                                                                                                                 �$POIO_GRP 1��������             �$POS_EDIT ��������                               �$POWERFL            �    �$PRGADJ ��������A�  A�  A�  ?   ?   ?      d    �$PRGNS_CFG ��������?�             @   <@�             %�                                                            �$PRGNS_GRP 2�������� �  \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                     �$PRGNS_PREF ��������      
    �$PRIORITY         ��   ��$PRMPDSPON            �    �$PRMPDSPOUT        �   �    �$PRODUCT_ID �������                       �$PROGGRP_TGL      ����    �$PROTOENT 1��������  (!AF_INET                              !tcp                                  !udp                                  !icmp                                 �$PROXY_CFG ��������  �    )� ****************************************   �)� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** �$PRO_CFG ��������    %�                                                          ?6�        ****/**/**/ **:**:**      %�                                         �                        A�    ,  �                                                                                     �$PRO_PREF ��������      
      �$PRPORT_NUM        �   �$PR_CARTREP  �������    �$PSKSTAT         �    �$PSSAVE ��������	2600H613                                              !�                                  !�                                  �                  	�          �        �                         �                      e�                                                                                                      �              !�                                  �$PSSAVE_GRP 1��������    �)                  ���������������������$PS_CONFIG ��������                     
          �  �   �2w��$PS_CP_CFG 2��������                                                         �$PS_CP_GRP 2�������   �         t�?g8���/[=
�?�?�  �^_7�þ7��H?��
�<�>TE}{tD*�    8���/[=
�?�?�  �^_7�þ7��H?��
�<�>TE}{tD*�        8�?�              ?�              ?�                  q8 $D    ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������       �$PS_MOTION 2�������� 
�                                %�                                      %�                                                                                                                  8�?�              ?�              ?�                                                                                                                                                                                                                                                                                                                             ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                    4%�                                   �A���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   '��%�                                     ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                     %�                                      ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   2 �%�                                   ����������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                     %�                                   EAL��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   '"%�                                     ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �[�%�                                   ����������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   U
�%�                                   � ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                      %�                                      ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$PURGE_ENBL         �   �$PWFENBDO            �    �$PWF_IO        �   �$PWRUP_DELAY ��������       �$PWR_HOT %������   �%�                                      �$PWR_NORMAL %�������%�                                      �$PWR_SEMI %�������%�                                      �$QSKIP_GRP 1��������  x 	                                      	                                                                              	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ����������������������������������������������������������$RBTIF      ����    �$RCVTMOUT        ��  ��$RDCR_GRP 1������� � 	 ?̏    E��UA�ҋC荽                 	 ��"9ŗ�            ����             	                                      	 ;��;QaT;\��;��;�	�<$D                    	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                   �$RDIO_TYPE  �������                                  �$REFPOS1 1�������� 
 x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS2 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS3 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS4 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS5 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS6 1��������  x�                                  	                                      	                                         �$REFPOS7 1��������  x�                                  	                                      	                                         �$REFPOS8 1��������  x�                                  	                                      	                                         �$REFPOSMASK 1��������     
   
   
   
   
   
   
   
�$REFPOSMAXNO  �������     
                     �$REMOTE  �������   �$REMOTE_CFG ��������          �$REPL_RANGE      ����   �$REPOWER ��������    �$RESM_DRYPRG %�������%�                                      �$RESTART ��������            �$RESUME_PROG %�������%�                                      �$RE_EXEC_ENB         �   �$RGSPD_PREXE         �    �$RGTDB_PREXE         �    �$RGTRM_PREXE         �    �$RMT_MASTER  �������    �$ROBOT_ISOLC  �������                 �$ROBOT_NAME �������KJLTVR411670R01       L T �$ROB_ORD_NUM ?�������  H613 �H895 �H895 \H895 P    �            ���     8�$RPC_TIMEOUT      ����   x�$RS232_CFG 1��������  LTEACH PENDANT                                  �                  Maintenance Conso                          "   �                  	Unbenutzt                                      �                  	Unbenutzt                                      �                  �$RS232_NPORT        �   �$RSCH_LOG ��������       		RSCH          �$RSMAVAILNUM        ��   �$RSPACE1 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                    ���������  ����������                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE2 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE3 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE4 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE5 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE6 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE7 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE8 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACEG ��������                           
 
                                                                                  ������������������������������������������������������������                                                                                                              d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������  `                  @   @   @                                                                           �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                ����������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  ��������������������� 
                                         �$RSPACE_MODE  �������    �$RSPACE_S ��������                                                                                                                          	                                     �$RSPCWORK_AD  �������~��$RSR  �������                  �$RSR_INTVAL        ��    �$RSR_OPTION         �   �$RTCFG ��������                      ?          �  �   �$RV_DATA_GRP 2�������   � D  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SAF_DO_PULS  ����   �������$SCAN_TIME        ��   �$SCR ����8

      
      
               
                                                                                                                                                                                                                                                                             �         2   2   
   
   d   
   d   2   d                        @                                                                          
                               P       
�� @B     T                                                                                    T D��                                                                                                                                                                                                                                                                                                                                                            @                    




                                             @         ;�o             p              
�t� �Di                        �                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                  �                                  0    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                                                                                                                                                                                                  �            �  �  � � � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �                   T                                                                                                                                                                                                                                                                                                                                                      �                                                       ��                                     	12345678    `!B  �            T                                                                                      T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T BH                                                                                                                                                                                                                                                                                                                                               T ;�j                                                                                                                                                                                                                                                                                                                                             T D�                                                                                                                                                                                                                                                                                                                                               T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   CH  A�               �          2                   
   d   
  �  	�     2                                                                                                       p  �                                  �                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                                                                                                                                                                                                                                                                                                                                                     �$SCR_GRP 1��� t �            	   � 	   � 	                                  	                                	                         @�          �      D�` D�@                 �    �                            R-2000iB/185L 567890  	R-2000iB  	R85L 678      
V06.10         	          
   
   
   
           	          �       �              	     	          � 	                                                                                                             ��H� 	     	   ��      OY]æ|XE�V�D�kB� :�.>C3�� 	 B�����:�@���8A �:�DE@                 <�Hæ}*E�V}D  	                                                            	                                         	                                     	 B���B�ffB�33B�  B�  B�  B�  B�  B�   	 A   A   A   A   A   A   @   @   @    	 @�  @�  @�  @�  @�  @�  ?�  ?�  ?�   	 BH  BH  BH  BH  BH  BH  A   A   A    	 F@ F�` F�`                          	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                            
                                         ?�  @�  @{f6                         	 @�  @�  @�  @�  @�  @�  @�  B�  B�  12345678901234567890                                                  A�                	                    	                                                                                                                                           P P P ( ( (                                                        �           	 	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	                                                              	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	                                                              	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	                                                              	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �$SEL_DEFAULT        ���   �$SEMIPOWERFL         �   �$SEMIPWFDO         �    �$SERVENT 1�������  L!DUM_EIP                             �j!AF_INET                           !FTP                                  !AF_INET                           !�                                    �!AF_INET                           !RPC_MAIN                            �!AF_INET                           !RPC_VISN                            �!AF_INET                           !TP_INPUT                            �d!AF_INET                           !
PMON_PROXY                          �e!AF_INET                           !TP_PROXY                            �f!AF_INET                           !RDM_SRV                             �g!AF_INET                           !R90                                 �h!AF_INET                           !
RPCM_PROXY                          �i!AF_INET                           !RLSYNC                              8!AF_INET                           !ROSIP                               �4!AF_INET                           !
CETP_MTCOM                          �k!AF_INET                           !	CETP_CONS                           �l!AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           �$SERVICE_KL ?%������  (%SVCPRG1                               %SVCPRG2                               %SVCPRG3                               %SVCPRG4                               %SVCPRG5                               %SVCPRG6                               %SVCPRG7                               %SVCPRG8                               %SVCPRG9                               %SVCPRG10                              %SVCPRG11                              %SVCPRG12                              %SVCPRG13                              %SVCPRG14                              %SVCPRG15                              %SVCPRG16                              %SVCPRG17                              %SVCPRG18                              %SVCPRG19                              %SVCPRG20                              %SVCPRG21                              %SVCPRG22                              %SVCPRG23                              %SVCPRG24                              %SVCPRG25                              %SVCPRG26                              %SVCPRG27                              %SVCPRG28                              %SVCPRG29                              %SVCPRG30                              �$SERVICE_PRG ?%������  (%                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       �$SERV_DEV �������MC:           �>��$SERV_MAIL      ����    �$SERV_OUTPUT      ����    �$SERV_REC 1�������   �    | 	   c  �  }  �  �  �   �         	                                  	    U      A            x         	                         Y         
 �X�[�6    	   2  t     *  �      ������ 	      �  �      6   �    ������ 	    b   ��������   �   �������� 	    ����   ��������L  �����������X��a6 2     	   �  s   �   �   �   �  ������� 	    n    �       I      %������ 	    ���������            $������� 	 ���f���F   ]�������A��������������X��6 2    	       �   �              ������ 	    �   �  a   p   t  
X   ������ 	 ���y   i����   �   �   ���������� 	 ����  d���)  �  ����  �������X��6    	   �     �      o      ������ 	       �          �      ������ 	    ���������            А������ 	 ��������      .���   C   ������X�6    	   g  �   �  
�  �  �    ������ 	       R   �   �   �       ������ 	    v   V�������<   n    �q������ 	 ��������  !������������   7������X�B@6 2     	    *  �     _      �    ������ 	       �  �   3      $   5������ 	 ���y   h����   �   �   ���������� 	 ����   ����  �  �����  4������X�+6 2     	    (  �     `      �    ������ 	       �  �   8      W   %������ 	 ���y   h����   �   �   ���������� 	 ����   ����  �  ����V  �������X�tC6    	   [  j     �  m  9    ������ 	    E  �        1   A    ������ 	    o   (��������   �   �������� 	 ����   1���#���$����  (����������X�xj6    	   ]  �   �  
Y  ~  �    ������ 	        y   �      �       ������ 	    v   V�������?   o    �q������ 	 ��������  �����������   3������X���6 2     	    &  �     _      �    ������ 	    
   �  
   5      B   >������ 	 ���y   h����   �   �   ���������� 	 ����   �����  m  ���
  [������    
 �Uv0�6 2     	                           ������ 	       �  �       �      ������� 	    ���������            ������� 	    P  ������������   ;  %|������U�=�6 2     	                           ������ 	       �  o       �       ������ 	    ���������            ������� 	    O   -   �������'   9  $�������X�;R6 2     	   �  H  �    �    ������ 	     �   �     "  �  
������� 	       &��������   i   � u������� 	 ����   �  U��������  �  !������Of*6    	   #  n  �  �  �  �  =������ 	       G  �       &   *    ������ 	    �������������   /     ������� 	    �   l  �����  �  #  �������X�hA6 2     	   �  V  �  �  �    )������ 	    �  �   �         	������� 	       &��������   i   � u������� 	 ����   �   ���������    i������Pq@�6 2     	                          ;������ 	       M  �       4      ������ 	    ���������            L������� 	    ����   �   ,����   5���P������P�e6 2     	                          ;������ 	       o  �       (      ������� 	    ���������            L������� 	    ��������   ���   ���{������Q1;�6 2     	                          C������ 	       y  �       "      ������� 	    ���������            L������� 	     �������   ���   ����������P��6 2     	                         A������ 	       �  �       *     	������ 	    ���������            L������� 	    ����  L   1����   J����������R8��6 2     	    
                     >������ 	       e         H      ������ 	    ���������            L������� 	 ��������   �   6���f   9����������     	                                      	                                      	                                      	                                      
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     	                                      	                                      	                                      	                                      
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     	                                      	                                      	                                      	                                      
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_RV 1�������   �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_TOP10 1�������   � 
 6T   6   _6    6 2  �6 .   6 i   6�   6 *   
6    76 s   �$SERV_TYPE      ����    �$SHELL_CFG ��������                                                                %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                                       �  �   %                                                                                                     �         �   2   d                                �$SHELL_CHK 1��������                                                                                                                                                                                                                                                                                                                                                                                  �$SHELL_COMM ��������                        �$SHFTOV_ENB         �    �$SHOW_REG_UI         �    �$SIMWAITENB            �    �$SIMWAITOUT        �   �    �$SIMWAITTIM       ��   �    �$SIMWAITVAL            �    �$SI_UNIT_ENB         �   �$SLC_RETRY         �   �$SMB_HDDN 2��������    ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  �������������������������$SMON_ALIAS ?e������ ( he�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      �$SMON_DEFPRO ������ *SYSTEM*    ��$SMON_RECALL ?}������ ( �}�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              �$SNPX_ASG 1�������� P 0 '%R[1]@1.1                              ?�      %                                    0?�      %                                     �?�      %                                    ?Z??�      %                                    �O�?�      %                                    o�o?�      %                                    �"?�      %                                    ���?�      %                                    � L?�      %                                    ���?�      %                                    �v�?�      %                                    ?�      %                                    �?�      %                                    ,?>?�      %                                    �O ?�      %                                    oho?�      %                                    �?�      %                                    ���?�      %                                    �0?�      %                                     ��?�      %                                    �Z�?�      %                                    ���?�      %                                    �?�      %                                    ?"?�      %                                    O�O?�      %                                    o L?�      %                                    ��?�      %                                    �v�?�      %                                    �?�      %                                    Ϡ�?�      %                                       ?�      %                                      �?�      %                                     c?�      %                                    :" ?�      %                                    ���?�      %                                    pP?�      %                                    ��?�      %                                    ���?�      %                                    �1?�      %                                    /K/?�      %                                    !�?�      %                                     �?�      %                                    /?�      %                                    -Q?�      %                                    
�c?�      %                                    Z?�      %                                     �b?�      %                                    <��?�      %                                    �x�?�      %                                    � �?�      %                                    � ?�      %                                    �l�?�      %                                    ��
?�      %                                    �?�      %                                    ?*?�      %                                     �O?�      %                                    oTo?�      %                                    ��?�      %                                    :�L?�      %                                    ޳?�      %                                    ��?�      %                                    ߂�?�      %                                    � ?�      %                                    � ?�      %                                    /J/?�      %                                    �?�?�      %                                    _t_?�      %                                     ?�      %                                     ��?�      %                                    �<�?�      %                                    ȿ�?�      %                                    �f�?�      %                                    ��?�      %                                    �?�      %                                    / .?�      %                                    �?�?�      %                                       ?�      %                                    ��l?�      %                                     %h?�      %                                      ?�  �$SNPX_PARAM ��������  �	�             P                           ��$SOFT_KB_CFG        ���    �$SOPIN_SIM  �������                                                  �$SRVQSTP_DSB  �������                                  �$SSR ������� � & FOLGE125 .......................0002        �$STHI_CHANGE         �    �$STHI_GRPNUM         �    �$STOP_ON_ERR         �    �$STOP_PTN ������C �$STRING_PRM         �   �$SVDT_GRP 1�������    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                   �$SVPRG_COUNT        ��    �$SVPRG_ENB         �    �$SVPRM_ENB         �    �$SVPRM_UPD 1������� T  
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                     �$SV_CTRL_NUM        
�   �$SV_GUN_CTRL 2��������                          
                        
                        
                           
                           
�$SYSDEBUG  ����   d�    �$SYSDSP_PASS       B?�    �$SYSLOG ��������         �^��                      �       UD1:\SYSLOG               �$SYSLOG_MPC ��������                                    �       UD1:\SYSLOG2              �$SYSLOG_SAV ��������                     UD1:\SYSLOGSV         �$SYSTEM_TIME 1��������  ( @�     .?V         #M$           �     @�     .C�         #M           �     @�     .C�         #M           �     @�     .C�         #M           �    �$T1SVGUNSPD        '�   ��$TASK_OPTION  ������   �   �$TA_DISP_ENB         �    �$TBCCFG ��������                                                 `                             	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                                                                	                                      	                                      	                                         ��������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������    �$TBCSG_GRP 2��������  �     
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ��� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������A��*SYSTEM*   V8.2306       4/24/2014 A t  *SYSTEM* *SYSTEM*  F�TBCPARAM_T   �$MC_MAX_TRQ  $MAX_TRQ_MGN  $MC_GRAV_MGN  $MC_STAL_MGN  $MC_BRK_MGN  $MC_NOLD_MGN  $SHORTMO_LIM  $SHORTMO_MGN  $MC_NOLD_TRQ  $J_LIN  $SPL1  $SPL2  $SPL3  $SPL4  $SPL5  $SPL6  $SPL7  $SPL8   8�TBC_GRP_T � $TBC_ACCEL1  $TBC_ACCEL2  $TBC_PATH1  $TBC_PATH2  $PATH_RATIO  $TBC_PARAM 2  	$CNT_SCALE  $SHORTMO_SCL  $MIN_ACC_UCA  $MIN_CAT_UMA  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2L_UPR_ANG  $J2L_LWR_ANG  $J2L_UPR_MGN  $J2L_LWR_MGN  $R_F2LSHRT  $R_F2LLONG  $MIN_F2LSHRT  $MIN_F2LLONG  $MIN_ACRL_S  $MIN_ACRL_L  $MIN_PAYLOAD  $HVAL   $HMGN   $FLEXL   ��TBJ_ACC_T  :$ACC_LEN1  $ACC_LEN2  $DEC_LEN1  $DEC_LEN2  $ACCEL_RATIO  $DECEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $F1DEC_I  $F2DEC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$DECTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT_ACC   	$J_STAT_DEC   	$M_STAT_ACC  $M_STAT_DEC  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $DEC2_STP   $AT_MODE  $AT_AXS   	$AC_ACC   	$AC_DEC   	$JK_ACC   	$JK_DEC   	$VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AA1  $AA2  $AA3  $AA4  $AA5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM  ���TBJCFG_T  � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $UPDATE_TIME  $TBJ_SELECT  $TBJ_STAT   $TJ 2 $JERK_CTRL  $MOTN_INF  $TBJ_DEBUG  $HAND_VB   �TBJOP_GRP_T  $ $F2MGN  $MINF2  $COMP_SW   ��TBPARAM_T � $$MR_MAX_TRQ  $MR_STAL_TRQ  $MR_BRK_TRQ  $MR_BRK_VEL  $MR_NOLD_VEL  $MA_LOAD_TRQ  $MD_LOAD_TRQ  $MAX_TRQ_MGN  $MA_GRAV_MGN  $MA_STAL_MGN  $MA_BRK_MGN  $MA_NOLD_MGN  $MD_GRAV_MGN  $MD_STAL_MGN  $MD_BRK_MGN  $MD_NOLD_MGN  $PTH_GRV_MGN  $PTH_STL_MGN  $PTH_BRK_MGN  $PTH_NLD_MGN  $DYN_FRC_MGN  $MR_NOLD_TRQ  $R_ACC_MGN  $R_DEC_MGN  $R_LONG_MGN  $J_ACC  $J_DEC  $DT_MGN  $SP1  $SP2  $SP3  $SP4  $SP5  $SP6  $SP7  $SP8  ��TBJ_GRP_T   $$TBJ_ACCEL1   	$TBJ_ACCEL2   	$ASYM_PARAM   $TB_PARAM 2 	$SHORTMO_SCL  $LONGMO_SCL  $MIN_ACC_SHM  $MIN_ACC_UMA  $SHORTMO_MGN  $LONGMO_MGN  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2J_UPR_ANG  $J2J_LWR_ANG  $J2J_UPR_MGN  $J2J_LWR_MGN  $INERTIA_VIB   $INERTIA_VI2   $IV_UNIT  $IV_UNIT2  $R_F2JACC  $R_F2JDEC  $R_F2JLONG  $MIN_F2JACC  $MIN_F2JDEC  $MIN_F2JLONG  $MIN_ACRJ_S  $MIN_ACRJ_L  $MIN_PAYLOAD  $HVAL   $HMGN   $HAXS   $FLEX    ��TCPPIR_T    $ENABLE_TCPP  $TCDELAY    ��TCPPSPEED_T  X $TCDELAY_MON  $VSPEED  $SPEED  $ACCEL  $TIMESTAMP  $PROG_SPEED  $MOTYPE  �TCPP_CFG_T 	 | $NUM_TCPPSEG  $GROUP_NUM  $TCPP_TIME  $WARNING_ENB  $OTF_TIM_ENB  $DEBUG_TASK  $DEBUG_MAIN  $TCPP_CMP_SW  ��TCPSPDCFG_T 
 � $TCDELAY  $HEARTBEAT  $SETUP_CFG  $SPD_MARGIN  $DEBUGFLG1  $DEBUGFLG2  $SPARE_STR1 $SPARE_STR2 $SPARE_LONG1  $SPARE_LONG2  $SPARE_REAL1  $SPARE_REAL2  `�TCPSPDOUT_T  p $ENABLE  $TARGET_TYPE  $TARGET_IDX  $MIN_VALUE  $MAX_VALUE  $MIN_SPEED  $MAX_SPEED  $GROUP_NO  �TP_THR_TABLE  $ $THR_ENB  $DI_NO  $DO_NO   ��THR_CFG_T  0 $MAX_IO_SCAN  $MIN_SCAN_TI  $SCAN_TIME  ��TIMER_T  � $COMMENT $TIMER_VAL  $STR_EPT_IDX  $STR_LIN_NUM  $END_EPT_IDX  $END_LIN_NUM  $TID_NUM  $DUMMY13  $PS_OVERFLOW   $OVERFLOW  $FLAG_TYPE  $FLAG_IDX  $GLB_TMR_ENB  $GLB_TMR_STR  t�TORQCTRL_T  X $DEBUG  $GRP_STT   $SBR_PAM21_V   T$SV_ERR_MOD   $SV_ERR_CLR   $ACTION  �TPGL_VIEW_T  4 $X  $Y  $Z  $WZ  $P  $R  $CAMERA    ��TPGL_UVIEW_T   $NAME $GIF }$VIEW D�TPGL_CAM_T  L $NAME $ID }$FID E$GIF }$NEARPLANE  $FARPLANE  $DISTANCE   �JOG_RAD_T   $JOINTS   	��TPGL_MSET_T    $NAME E$ID }$TIMECONST  ��TPGL_CONF_T � $MOUNT ?� $LOCK_FOLLOW  $DBGLVL  $GLDBGLVL  $TEST_XML }$TEMPINT   $TEMPSTR ?� $USER_VIEWS 2 $CAMERAS 2 $TEMP_LOCS 2 $SCENE_VIEW 2  $KAREL_TMO  $TPDRAW_TMO  $JOG_VECLEN  $JOG_RADIUS 2 $CHECK_TOOLS  $CHECK_VIS  $REG_VIS32  $REG_VIS64  $MACHSET 2 $CONT_IDX  $DUMMY29  $VISIBLE   @$RAIL_BOXES   $ROBOT_XML ?� $SHOWWARN   $PS_CONTROLM   $CONTROLMAX  $CONTROLMASK   $FP_TO_FK ! �TPGLMACH_T   $JOINTS   	 ��RECLOC_T   $SLOTS !   ��TPGL_OUT_T  X $VIEWS 2 $SELECTED ?� $PIP_XML }$NODEVIS   @$MACHINES 2 $RECORDEDLOC 2 H�TPP_MON_T  D $GLOBAL_MT  $LOCAL_MT  $MON_NUM  $GMON_TID  $SYSMON_ADR  �TPSTRTCHK_T  , $ENABLE  $ALLOW_NAME $ALLOW_LINE   ��TPVWVAR_T  � $TPVIEW_ENB  $PREV_RTN  $EDIT_RTN  $VSHWRK  $DEBUG  $DISPLAY  $INDENT1  $INDENT2  $HEAD1 $HEAD2 $EDIT_KEY  $TCPSPD_KEY  $JMPCALL_ENB  @�TRACE_CFG_T  D $ENABLE  $ITEMS  $CHANNELS  $DEBUG  $TICKS  $MIN_MM  �TRACE_CHNL_T  @ $ITEM_NUM  $TCP_GP_NUM  $VISIBLE  $STYLE  $COLOR    ��TRACE_ITEM_T  t 
$PRG_NAME %$VAR_NAME =$DESC !$UNITS $TYPE  $IO_TYPE  $PORT_NUM  $SQUARE  $SLOPE  $INTERCEPT  ��TSCFG_T  $GRP_MASK  $MODE_MASK  $STATUS  $OPT_VAL  $SIZE  $FNAME_TYPE  $PS_PROC   $PROC  $OUTPUT  $OUTPUT_DONE  $AXS_MSK_ENB  $AXIS_MASK   $CUR_RECTIME  $TOT_CHN_NUM  $MINFREQ_US  $SETFREQ_POW  $LPARAM   
$FPARAM   
$PATH_NAM $DUMMY19  $DUMMY20   ��TSR_GRP_T  l $MR_MAX_TRQ   	$MR_STAL_TRQ   	$MR_BRK_TRQ   	$MR_BRK_VEL   	$MR_NOLD_VEL   	$MA_LOAD_TRQ   	$MD_LOAD_TRQ   	$MA_GRAV_MGN   	$MA_STAL_MGN   	$MA_BRK_MGN   	$MD_GRAV_MGN   	$MD_STAL_MGN   	$MD_BRK_MGN   	$MJ_ACC_MGN   	$MC_ACC_MGN   	$MC_STAL_MGN   	$MC_BRK_MGN   	$MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	��TSSCB_T ! h $DSP_NO  $DSPAX_NO  $DATA_SEL  $OUT_CHANNEL  $ADDRESS  $BIT_SHIFT  $USE_2CH  $MONITOR  �TXSCREEN_T " $ $DESTINATION }$SCREEN_NAME �&��REQ_DATA_T # T $ERR_TYPE  $ERR_GRP  $ERR_AXIS  $AXIS_TYPE  $ERROR_DIST  $ERR_TIME   ��UECFG_T $ � 	$CHK_VERSION  $RSM_CHK_ENB  $UNEXCEP_ENB  $RSM_THRS_R  $RSM_THRS_L  $UNEX_THRS_R  $UNEX_THRS_L  $REQ_COUNT  $REQ_DATA 1# 
�UEGRP_T % 0 $ERR_COUNT  $PROGMTN_FLG  $CURR_POS   	��UI_MENHIS_T & 8 $HIST_HEAD  $HIST_ENTRY ?� $DUMMY2  $DUMMY3  8�UI_MOUSE_T ' @ $ACTION  $BUTTON  $ROW  $COLUMN  $TIME  $RESERVED  �UI_PANEDAT_T ( � $PAGEURL }$FRAME )$HELPURL }$PARAMETER1 )$PARAMETER2 )$PARAMETER3 )$PARAMETER4 )$PARAMETER5 )$PARAMETER6 )$PARAMETER7 )$PARAMETER8 )$INTERVAL  $PANESTATE  $DUMMY14  $MOUSE '�UI_USRVIEW_T ) < $MENU $CONFIG $FOCUS $PRIM m$DUAL m$TRIPLE m�UNDO_CFG_T *  $UNDO_ENB  $WARN_ENB  ��USER_INFO_T + 8 $USR_PROG %$TASK_ID  $USR_POSIDX  $USR_PR_USE  �USER_TOOL_T , 4 $X  $Y  $Z  $W  $P  $R  $TOOL_NUM  ��USER_UFRAM_T - 4 $X  $Y  $Z  $W  $P  $R  $UFRAME_NUM  �USER_OFFST_T . D $TOOL_OFST 1, $UFRAME_OFST 1- $GUN_WIDTH   $ENB_SUBNUM   
�USRTOL_GRP_T / @ $DIST_TOL  $ORNT_TOL  $RAUX_TOL  $TAUX_TOL  $ENABLE  �VCCM_CFG_T 0  $SC36MFB1ENB   4�VCMR_CAM_T 1h $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DETECT_TYPE  $DRIVE_TYPE  $SET_VTCP  $DEBUG_CODE  $DMY_UBYTE  $CAMERA_NAME %$DISTORTION1  $DISTORTION2  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $HANDEYE  $EXPOS_TIME  $NUM_MUL_EXP  $FOCAL_DIST  $GD_SPACING  $TRGT_DIST  $TRGT_W  $TRGT_P  $TRGT_R  $NUM_RETRY  $UTOOL   t�VCMR_TRGT_T 2  $TARGET_PNT   x�VCMR_CRPR_T 3 d $AXIS_FLAG   	$NUM_AXS_REP  $SWING_ANG   $NUM_MS_POSE  $BASE_POSE   	$EVALUE_IDX   `�VCMR_CHKM_T 4 @ $EVALUE_IDX  $MAX_MS_ERR  $MEAN_MS_ERR  $WORST_POSE   ��VCMR_MRCV_T 5 � $ORG_MST_CT   	$ORG_UFRAME   $ORG_REF_POS   	$ORG_REF_CT   	$RCV_ANG_PAM   	$NEW_MST_CT   	$NEW_UFRAME   $NEW_REF_POS   	$NEW_REF_CT   	$EVALUE_IDX  $MAX_RC_ERR  $MEAN_RC_ERR  $WORST_POSE  $MASTER_TIME  $DEBUG_MODE   ��VCMR_GRP_T 6 � $STAT_FLAGS  $MENU_CODE  $GROUP_NUM  $UTOOL_NUM  $CAMERA 1$TARGET_ID 22 $CREATE_PRG 3$DATA_ID  $CHK_RESULT 4$RECOVERY 5$EXT_INT1  $EXT_INT2  $EXT_INT3  $EXT_INT4  $EXT_REAL1  $EXT_REAL2  $EXT_REAL3  $EXT_REAL4  �VISION_CFG_T 70 &$DATA_PATH  $DATA_CACHE  $LOG_PATH  $LOG_EXPATH  $LOG_TIMEOUT  $MC_LIMIT  $FR_LIMIT  $TD_LIMIT  $DEBUG_MODE  $HOST_NAME  $COMM_PORT  $ROBOT_NAME  $FLAGS  $MAX_PAGES  $MIN_VPOOL  $VPOOL_SZ32  $VPOOL_SZ64  $VPOOL_SZ128  $VPOOL_SZCAL  $VPOOL_LIM  $VPOOL_WAIT  $TMPPOOL_LIM  $FAILIMG_IDX  $LOADIMG_IDX  $NUM_IMREGS  $IMREG_SIZE  $GPM_CANDMAX  $NUM_ASYNBUF  $NUM_VRTDBUF  $VRTDBUF_SIZ  $TOLE_2D_Z  $TOLE_2D_WP  $PC_SETUP  $LOGQUE_MAX  $ECCU_RETRY  $VEMT_PATH  $VEMT_LIMIT  $VIRCIMG_SIZ  T�VISION_GRP_T 8  $BACKLASH   	�VLEXE_CFG_T 9 D $ENABLED  $DATE  $FLDR_INDEX  $FILE_INDEX  $REC_INDEX  |�CUSTOMMENU_T : $ $TITLE $PROG_NAME %$OPTION  �VSHIFT_CFG_T ;` $DATA_NAME 	$CAMERA_NAME %$EXPOSURE  $WIN_RADIUS  $WIN_POS_X  $WIN_POS_Y  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $LIM_DIST  $LIM_ANGLE  $LIM_TILT  $LIM_SCORE  $LIM_CNTRST  $WARN_DIST  $WARN_ANGLE  $WARN_TILT  $WARN_SCORE  $WARN_CNTRST  $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DUMMY23  $USED_CAMTYP    �VSMO_CFG_T <  $ENABLE  $ADJUST_TIME  �WAIT_DATA_T =  $PROG_NAME %$LINE_NUM  �WV_AXSRST_T >   $AXIS_MASK  $THRESHOLD   ��ZABC_GRP_T ?  $ZABC_MODE   
 ��ZMPCF_GRP_T @   $ZMP_ENB  $ZMP_DMY_LNK   
��ZMPOS_GRP_T A � $M_POS_ENB  $CMCMD_SCL  $CART_MCMD   	$P_ACT $J_ACT   	$P_DES $J_DES   	$P_DES2 $J_DES2   	$UXWPR_ENB  $UXEUL_ENB  $UXWPR_ACT   $UXWPR_DES   $UXEUL_ACT   $UXEUL_DES     ��ZP_CFG_T B  $ENABLE  $DEBUG   ��ZP_CYLINDER_ C 8 $RADIUS  $HEIGHT  $PROG_NAME ?( $LINE_NUM   D�ZP_GRP_T D � $OPTIONS   
$BREAK_TIME  $WORK_SHIFT  $ENABLE  $RV_LIFE   	$SHIFT_OVC   	$PART_ID  $OPTM_RATE   
$MAX_I_RATE  $MAX_DI_RATE  $TRACE_ENV  ��ZP_SPHERE_T E , $RADIUS  $PROG_NAME ?( $LINE_NUM   ��$TBC_GRP 2������� d � �?    	 HD)�?�  ?�  ?   ?   ?fff?�  ?�  C��nA�                                  D)�?�  ?�  ?   ?   ?fff?�  ?�  C��nAP                                  D)�?�  ?�  ?��?��?�  ?�  ?�  C��nA�                                  C?�  ?�  ?fff?fff?fff?�  ?�  CA�BP                                  C?�  ?�  ?fff?fff?fff?�  ?�  CA�BP                                  C?�  ?�  ?�  ?�  ?�  ?�  ?�  CA�BP                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  ?�  ?�     �  	V3.00     	r85l      	****      	�          B�                  ?L��?�33   x   �?�  ?�                                            ?���Cz                                          ������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  �������������������������������������$TBJCFG �������                 �                                     �                                                 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                              	                                      	                                      	                                      	                                      	                                                                                      	                                      	                                      	                                         ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������                                             �$TBJOP_GRP 2�������  ?���CH     	����������������������������$TBJ_GRP 2������� � 	 ����X�       	 �X^ �,X        @   ?�   	 �D)�D)�D)�C2
C랔        ?�  ?�  ?333?333?�  ?�  ?333?333?�  ?�  ?�  ?�  ?�  <^�%C��n?fff?�=q?L��A�  A@      ?�                              D)�D)�D)�C2
C래        ?�  ?�  ?333?333?�  ?�  ?333?333?�  ?�  ?�  ?�  ?�ff<�7�C��d?���?���?���A�  Ap      ?�                              D)�D)�D)�C2
C랔        ?�  ?�  ?333?333?�  ?�  ?333?333?�  ?�  ?�  ?�  ?�  <�\�C��n?�ff?Ǯ?�  B  A�      ?�                              CCCC���C�p�        ?�  ?�  ?fff?fff?fff?�  ?fff?fff?fff?�  ?�R?�R?L��;���CA�?���?���?�  B�  B                                      CCCC���C�p�        ?�  ?�  ?fff?fff?fff?�  ?fff?fff?fff?�  ?&ff?&ff?L��;YQ@CA�?fff?�=q>���B�  B                                      CCCC���C�p�        ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?L��?L��?�  <RxCA�?�33?�
=?�  B�  B                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      C�         �  0?�  ?�  	V3.00     	r85l      	****      	�          B�                    F�� F�� F�� G� G@ G;� GZ� Gz  G�� G� G�� G� G�x G�� H� HL H'� H7� HG8 HV�   F�� F�� F� F�0 G� G� G ( G3� GG8 G^� Gz  G�� G�@ G�� G�\ G�� G�` G�� H� HR =u=+?�  ?�  ?�     p   p   �?�  ?�                                                          ?�  @   ?�  ?�                               	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  �������������������������������������$TCPPACTSW  ������     �$TCPPIR �������   CH  �$TCPPSPEED ������ CH                      t�?�        �$TCPP_CFG 	�������                          �$TCP_SPD_CFG 
�������     �m   :�o        �              �                              �$TCP_SPD_NUM      ����   
�$TCP_SPD_OUT 2������� 
                                                                                                                                                                                                                                                                                                              �$TCZEROSPD              �$TESTPARS  ������   �    �$THRESTABLE 1�������                                                                                                 	           
                                                                      �$THRRDITABLE 1�������                                                                                          �$THRRDOTABLE 1�������                                                                                          �$THRSDITABLE 1�������                                                                                                                                                                                                                                                                                                                                                                                                   �$THRSITABLE 1�������                                                                                                             	           
                                                           �$THRTABLENUM  �������          �$THR_CFG �������   
   @   ��$TIMEBF_TTS         
�   �$TIMEBF_VER        
�   �$TIMER 1�������   8�                   �
� 
�  ��         �       �                   �
� 
�  ��         �       �                    7�
� 
�  ��         �       �                  ����� ��  H��        �      �                    �@� 8  ��         �       �                    �p	J 	S  ��         �       �                  �A�c���  H��         �      �                  �*c���  H��         �      �                  �C�c���  H��         �      �                   ��@� ��  H��         �      �               ���    �  �   ��         �       �               ʿ������ 	��  H��        �      �                  OJ��� ��  H��         �      �                   	O< <  ��         �       �               �    �  �   ��         �       �               SSS    �  �   ��         �       �                �    �  �   ��         �       �                      �  �   ��         �       �               X     �  �   ��         �       �                      �  �   ��                   �                     �  �   ��                   �               kU    �  �   ��                   �               7     �  �   ��                   �               �O�    �  �   ��                   �               MR     �  �   ��                   �               N ?    �  �   ��                   �               � �    �  �   ��                   �               ���    �  �   ��                   �               ED     �  �   ��                   �               ���    �  �   ��                   �                �    �  �   ��                   �               L      �  �   ��                   �$TIMER_NUM        @�    �$TMI_CHAN          �    �$TMI_DBGLVL         �    �$TMI_ETHERAD ?�������  0000:e0:e4:34:0e:af 0000:e0:e4:34:0e:b0 �                  0000:e0:e4:34:0e:b2 �$TMI_ROUTER !�������!ROUTER                            �$TMI_SNMASK ?�������  255.255.255.0     255.255.255.0     255.255.255.0     255.255.255.0     �$TOOLOFS_DIS         �    �$TORQCTRL ������                                       T                                                                                                                                                                                                                                                                                                                                                                                                                         �$TPE_DETAIL         �   �$TPGL_CONFIG ������  �?/cell/$CID$/grp1              ?�                                                                                                  �/cell/$CID$/grp2                                                                                                                  �/cell/$CID$/grp3                                                                                                                  �/cell/$CID$/grp4                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                             }�                                                                                                                                                                                  ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                    �User View 1           }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345 ���������������������User View 2           }�                                                                                                                              ���������������������User View 3           }�                                                                                                                              ���������������������User View 4           }�                                                                                                                              ���������������������User View 5           }�                                                                                                                              ���������������������User View 6           }�                                                                                                                              ���������������������User View 7           }�                                                                                                                              ���������������������User View 8           }�                                                                                                                              ��������������������� lCamera 1              }�                                                                                                                              E�                                                                      }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345             Camera 2              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 3              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 4              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 5              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 6              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 7              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 8              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 9              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 10             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 11             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 12             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 13             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 14             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 15             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 16             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   
   (  �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������                 �E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ����� @ ����������������������������������������������������������������  ��������  ��)frh:\tpgl\robots\r2000ib\r2000ib_185l.xml                                                                                                                                                                                                                 � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                            ���������     ����������������  88�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  �$TPGL_OUTPUT ������   ���?�              ?�              ?�                  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     }�                                                                                                                               @ ����������������������������������������������������������������  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  �  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8�����������������������������������������$TPOFF_LIM      ����   �$TPON_SVOFF         �    �$TPP_MON �������          2        �$TPSTRTCHK �������    �                  �$TPVTCOMPAT         �    �$TPVWVAR �������                   �                  �                       �$TP_DEFPROG %�������%FOLGE125                              �$TP_DISPLAY  �������    �$TP_INST_MSK  �������          �$TP_INUSER         �   �$TP_LCKUSER         �    �$TP_QUICKMEN         �    �$TP_SCREEN �������t_sc  �$TP_USERSCRN �������t_sc  �$TP_USESTAT         �    �$TRACE_CFG ������         	       
?�  �$TRACE_CHNL 2������ 	                 �                 �                 �                 �                 �                 �                 �                 �                 � �$TRACE_ITEM 2������  �%$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          �$TSCFG ������                 �  �                                                   
                                          
                                         UD1:\               ���$TSR_GRP 1 ������ � 	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678  �$TSSCB 2!������                                                                                                                                                                                                  �$TX_SCREEN 1"������ 
 �}ipnl/pnlgen.htm                                                                                                               Panel setup               }	index.STM                                                                                                                     
Robot Info e              }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          �$UALRM_MSG ?������� 
  �                              �                              �                              �                              �                              �                              �                              �                              �                              �                              �$UALRM_SEV  ������� 
   �$UECFG $������           @�  A�  A   B�   N� 
   �          B�
�X�^V  �          B�7 X��a  �          BȲ�X�H�  �          B���X�PG  �          BȺpX�Q  �          BȾ�X�Q�  �          B�T�X�X�  �          B�İX�\�  �          B�@X�K�  �          B��@X�Z��$UEGRP 2%������  0 N�    	 ?�ٿ2��Vv����U>2��7�SE@                  	                                              	                                              	                                     �$UI_DEFPROG ?%�������  (%UP002 11                              %$UP222...........................0050  %�                                      %�                                      %�                                      %�                                      %�                                      %�                                      �$UI_INUSER  �������                                  �$UI_MENHIST 1&������  (   ��-/SOFTPART/GENLINK?current=editpage,FOLGE020,1 8 ...................0050,9                                                         �'/SOFTPART/GENLINK?current=menupage,18,1  11,3                                                                                     �-/SOFTPART/GENLINK?current=editpage,FOLGE125,2  ....................0050,9                                                         �'/SOFTPART/GENLINK?current=menupage,98,1 011,7                                                                                     �+/SOFTPART/GENLINK?current=editpage,UP002,27 1 .....................0050,8                                                         �)/SOFTPART/GENLINK?current=menupage,1110,1 6 1                                                                                     �'/SOFTPART/GENLINK?current=menupage,71,1 018,23                                                                                    �'/SOFTPART/GENLINK?current=menupage,37,1 020,1  ....................0050,8                                                         ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ���$UI_PANEDATA 1(������  	�}/frh/cgtp/doubdev1.stm 8981&action=100                                                                                        )prim                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ��    ��\    }/frh/cgtp/doubdev2.stm mode=1                                                                                                 )dual                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ��    B�����}  frh/cgtp/tdev3.stm                                                                                                           )  hird                                     }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �   	 Bi����}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}�                                                                                                                              )�                                          }�                                                                                                                              )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          ��������������$UI_POSTYPE  ������� 	                                     �$UI_QUICKMEN  �������                                  �$UI_RESTORE 1)������  ��                                             �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �$UI_SCREEN ?�������  u1sc  u2sc  u3sc  u4sc  u5sc  u6sc  u7sc  u8sc  �$UI_USERSCRN ?�������  u1ks  u2ks  u3ks  u4ks  u5ks  u6ks  u7ks  u8ks  �$UNDO_CFG *�������      �$UPDATE �������KS_24 �$USER_INFO 1+�������  0%  P022                                         %                                               %                                               %                                               %                                               %                                               %                                               %                                               �$USER_OFFSET .�������                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                                   
                                         �$USEUFRAME         �   �$USRTOL_ABRT         �    �$USRTOL_ENB         �   �$USRTOL_GRP 1/�������  Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz     Cz  A�  A�  Cz     Cz  A�  A�  Cz     �$USRTOL_MENU            �    �$USRTOL_MSK         �    �$USRTOL_NAME %�������%�                                      �$VCCM_CFG 0�������    �$VCMR_GRP 26������               	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                    �$VISIONTMOUT        ��  ��$VISION_CFG 7�]p�^� FR:\VISION\DATA\                   �� MC:\VISION\LOG\                    UD1:\VISION\EXLOG\                  ' B@ �� ��     �                                                                                  �  =	 1- n6  -��         B@         ,             =���=���            MC:\VISION\TRAIN\                       �$VISION_GRP 28������  ( 	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���            �$VLEXE_CFG 9������    1-e            �$VMPHASE  ������          �$VSHIFTMENU 1:������ 
 <�              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���	LIVE/SNAP     %vsflive                               ���VISION SETUP  %vsfmenu                               ����              %�                                      ����$VSHIFT_CFG ;�������	�          %�                                        �5   @   �  @����       A�  B8  B  B�  Ap  Ap  B  A�  B�  B    �  ���������$VSHIFT_MEP        ���   �$VSMO_CFG <������    �z  �$WAITDINEND        �   �    �$WAITDINOK            �    �$WAITDINOUT        �   �    �$WAITDINST        �   �    �$WAITDINTIM       ��   �    �$WAITGINEND        �   �    �$WAITGINOK            �    �$WAITGINOUT        �   �    �$WAITGINST        �   �    �$WAITGINTIM       ��   �    �$WAITRELEASE         �    �$WAITTMOUT        ��  ��$WAIT_ACTIVE         �    �$WAIT_DATA =�������%  OLGE125........................0001      �$WAIT_RDISP         �    �$WV_AXSRST 2>�������                                  �$WV_GRP_IR  ������ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �$ZABC_GRP 1?������  , 
        2                                 
        2                                 
        2                                 
        2                                �$ZMPCF_G 1@�������  0     
                                              
                                              
                                              
                                         �$ZMP_GRP 1A������  �      � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��  �$ZPCFG B�������        �$ZP_CYLINDER 2C�������  �          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZP_GRP 2D�������  � 
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�  �$ZP_SPHERE 2E�������  �      ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZZZ         ��    