A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DMR_GRP_T  � $MASTER_DONE  $OT_MINUS   	$OT_PLUS   	$MASTER_COUN   	$REF_DONE  $REF_POS   	$REF_COUNT   	$BCKLSH_SIGN   	$EACHMST_DON   	$SPC_COUNT   	$SPC_MOVE   	$ADAPT_INER   	$ADAPT_FRIC   	$ADAPT_COL_P   	$ADAPT_COL_M   	$ADAPT_GRAV   	$SPC_ST_HIST   	$DSP_ST_HIST   	$SHIFT_ERROR  $SPC_CNT_HIS   	$MCH_PLS_HIS   	$ARM_PARAM   d$MASTER_ANG  $DSP_ST_HIS2   	$CLDET_CNT   	$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$GRAV_MAST   P�FMS_GRP_T t *$REM_LIFE   	$NT_LIFE   	$T_LIFE   	$CLDET_ANG   	$CLDET_DSTB   	$NT_LIFE_0   	$T_LIFE_TEMP   	$REM_LIFE_0   	$GRP_CL_TIME  $PCCOMER_CNT   	$FB_COMP_CNT   	$CMAL_DETECT   	$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $DTY_STR_T  $DTY_END_T  $CLDET_CNT   	$CLACT1   $CLACT2   $CLACT3   $CLACT4   $CLACT5   $CLACT6   $CL_OVR   $CLOMEGA1   $CLOMEGA2   $CLOMEGA3   $CLOMEGA4   $CLOMEGA5   $CLOMEGA6   $CL_FRMZ   $CLDEPT_IDX   $CLCURLINE   $CLDEST1   $CLDEST2   $CLDEST3   $CLDEST4   $CLDEST5   $CLDEST6   $CLNAME ?( �PLCL_GRP_T  � 	$CALIB_STAT  $TRQ_MGN   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	��VCAX_REFA_T  @ $REF_FACTORY  $NUM_SET  $MAST_TO_REF  $PRE_MST2REF   <�VCAX_REFD_T  , $COMMENT $REF_UPDATE  $REF_AXIS 2 	L�VCAX_REFS_T  8 $STEP_MS_ENB  $NUM_SET  $STEP_DATA  $PRE_STEP  �VCAX_REFM_T   $IS_SET  $MASTER_COUN  �VCAX_REFG_T  0 $REF_DATA 2 
$REF_STEP 2 	$PRE_MASTER 2 	�$$CLASS  ������       �$DMR_GRP 1 ������      	                                      	                                      	  ��x? �?��')��w��,	r                 	                                      	                                      	                                    	                                	 �X^� ���LM���i�s(����             	                                      	                    	                    	                    	                    	 ���� �� )       	              	 B B    B                     	 ���������K�_�����.��             	  �����m���?�'��wV�,	5             d                                                                                 =L��                                    ?�                              @�                                                                                                                                                                                                                                                           	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 �����$FMS_GRP 1������  	 I*eG�[�H0e�H�S"I�V�I=Y             	 M�9O�N�-sJ�BI��QI�=             	 B�  B�  B�  B�  B�  B�               	 B���BO��'Bޜ!©>�A+��             	                                      	 N�^=P�q�P7D�L�7>K��bK:A              	 A��iA��iA��iA��iA��iA��i             	 I*�G�^H0f�H�S�I�WI=�            X�}� 	                                     	                                  	                                                                Wy<WyBX�}X�}�X�}�O���PJ^�PU�V�V�V�V�(Wx�Wx�Wx�Wx�WyWyWyWy(X��X�. 	    !                                �������� ��
�y�
���p�R��߳�p�*���Q�������)������!��,��o"��N���2���O������d  �<��Ia��n��P��4-?3�5�-��[��p����_4��6������X�����+v�9B   6�U 6�K��S���?:��O����!����������
{ 7r� 7j� 7L� 7.� 7� 6�� 6�" 6��  Cz�Cxl�u��r��n)�Ux'� }S�}Qa}N&}S�C��C��C�JC��C��C�C}�C{�  ��^@��^@������������s��L�s '�s��s�%�s���s����Y���Z���[Y��\"��]H��]���]���^  �?
��?�Iظ�I�<�I�>��a=�H7��`���lZ��l���m	��lU�?
m�?	�?	f�?	��?	��?
�?
b�?
�           d         d   d   d   
   
   
      
                                   ����  ����  �                                             ����  �����������|F��������   ����           ����                                ����     5|���  4�                          ����                   ����    �������5���%��ƃ      ������������        ����   ����                  ���5   �������o����������������       ����        ��������                    ����         4   @  �               ����    ����       ����             e   e   e   e   e   e   e   e   f   f   f   f   e   e   e   e   e   e   e   e                                                                                          �   N   N      M      D   D   D   C                          ?�E�?�L�?��E?�;+?�L�@s?�:_@s?���?��?� �?��V?��t?��S?�b?��?�)*?�3�?�>�?�B�  ?�\?��?�?�?ʺ>y~F?y�>y~C?`�?Z�?��?Q/?Q�?V�?a�?J~?pV?y�?��?yN  ��Ŀ�=��e����������]Կ�0��]�=ϴ�=��7=͟�=�hO���������������꿌�|��衿��2���  ?�~�?�}�?��d?���?��?[V�?��p?[Vҽ��s�������J����?ل�?ـ�?��?ـ7?ـ?�2?�z??ق�  ���Ͽ��¿�ĵ��Ŀ�j��8������8���cٿ�^Y��a$��_O�������7�������u������ڿ��(���o  ?��_?��>?�g>?�u>?�&@ �>?�w@ �@:�@<S@;@<D?���?��\?��9?���?��A?��y?��K?��o  ,($UP001                                     ($UP001                                     ($VW_USER                                   ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP021                                     ($UP021                                     ($UP021                                     ($UP021                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                     ($UP001                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      �$PLCL_GRP 1������� D    	 ?�  ?�  ?�  ?�  ?a��?w�?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$VCAX_REF_GR 2������ t 
 �REFERENCE 1        	                                                                                                                                                 REFERENCE 2        	                                                                                                                                                 REFERENCE 3        	                                                                                                                                                 REFERENCE 4        	                                                                                                                                                 REFERENCE 5        	                                                                                                                                                 REFERENCE 6        	                                                                                                                                                 REFERENCE 7        	                                                                                                                                                 REFERENCE 8        	                                                                                                                                                 REFERENCE 9        	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE2_1       	                                                                                                                                                 REFERENCE2_2       	                                                                                                                                                 REFERENCE2_3       	                                                                                                                                                 REFERENCE2_4       	                                                                                                                                                 REFERENCE2_5       	                                                                                                                                                 REFERENCE2_6       	                                                                                                                                                 REFERENCE2_7       	                                                                                                                                                 REFERENCE2_8       	                                                                                                                                                 REFERENCE2_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE3_1       	                                                                                                                                                 REFERENCE3_2       	                                                                                                                                                 REFERENCE3_3       	                                                                                                                                                 REFERENCE3_4       	                                                                                                                                                 REFERENCE3_5       	                                                                                                                                                 REFERENCE3_6       	                                                                                                                                                 REFERENCE3_7       	                                                                                                                                                 REFERENCE3_8       	                                                                                                                                                 REFERENCE3_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE4_1       	                                                                                                                                                 REFERENCE4_2       	                                                                                                                                                 REFERENCE4_3       	                                                                                                                                                 REFERENCE4_4       	                                                                                                                                                 REFERENCE4_5       	                                                                                                                                                 REFERENCE4_6       	                                                                                                                                                 REFERENCE4_7       	                                                                                                                                                 REFERENCE4_8       	                                                                                                                                                 REFERENCE4_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                         