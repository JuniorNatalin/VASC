A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DRYRUN_T   � $DRYRUN_ENB  $NUM_PORT  $NUM_SUB  $STATE  $TCOL_SYSPT  $PMC_SYSPT  $GRP_MASK  $STEP_MOTION  $LOG_INFO  $TCOL_SAVE  $FLTR_EMPTY  $PROD_START  $ESTOP_DSBL  $POW_RECOV  $OPR_DSBL  $SAW_PROG %$INIT_PROG %$RESUME_TYPE  D�DRYRUN_PORT_  4 $TYPE  $FST_IDX  $LST_IDX  $STATIC_PORT  ��MIX_BG_T  4 $PROG_NAME %$MODE  $STATUS  $MODIFY_TIME  ��MIX_MKR_T   $LINE   $LINE_SIZE   ��MIX_LOGIC_T , $USE_FLG  $USE_MKR  $USE_TCOL  $USE_TCOLSIM  $NUM_FLG  $NUM_MKR  $NUM_BG  $NUM_SCAN  $MAXNUM_SCAN  $MINNUM_SCAN  $ITEM_COUNT  $PROC_TIME  $MAX_TMR_VAL  $TCOL_LINE $TCOL_ENB  $TCOL_SIM  $TCOL_STAT  $SAVE_IDX  $SAVE_LINE $TCOL_WARN  $BG_HITEM  $INST_CHK  �$$CLASS  ������   5    5�$DRYRUN  ������5�      c                        ����                   %VAGSAW                                %VAGTPINI                                 �$DRYRUN_PORT 2������5� c    "      $             d                   )     �                                             	  	                    �  �         �  �         �  �         �  �         �  �                    !  8         c  c         h  i         l  l         y  �         �  �         �  �         �  �                      	                      2         9  ;         A  P         a  x         �  �         �  �         �  �         �  �         �  �         �  �         �  �         �  �           !         )  +         C  C         H  I         L  L         Q  q         y  {         �  �         �  �         �  �         �  �         �  �         �  �         �  �         	  	         !  3         7  7         I  I         a  s         w  w         �  �         �  �         �  �                                 1  A         V  a         v  �       )   D   G       )   M   P       )   y   z       )             )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )           )  !  !       )  2  2       )  J  J       )  A  A       )  P  P       )  `  c       )  e  e       )  u  x       )  z  z       )  �  �       )  
  9       )  �  �       )  �  �                                                                                                    �$DRYRUN_SUB ?������5�  FOLGE         UP         0  MAKRO         SUCHL         BIN1        D�$MIX_BG 2������5�  4%MAKROSP1                                    J{��%MAKROSP2                           </t      J{��%MAKROSP3                           h=3      ����%MAKROSP4                           5-1      ����%MAKROSP5                           ="4      ����%MAKROSP6                                    ����%MAKROSP7                           ame      ����%MAKROSP8                            �      J{���$MIX_LOGIC ������5�                  �              X  ����   2tq* _t
 Pq* _t* q* _t                                                                                                                                                                                                                                               ����  s2tq* _t
 Pq* _t* q* _tBqu) Hqu) Iqs) Zr) \ttq�tt�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������              �$MIX_MKR 2������5 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ds
 q
 q
t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   _ds
�qu
�q
�q
�qssu
�q
�tr�tqu
qu
q�t                                                                                                                                                                                                        `ds
Jqu
Lqu
Kq
Mqu�qs)Arskq) �trsq) �ttt                                                                                                                                                                                                       adss
�q�r)8tq
BqBqu) Hqu) Iqs) Zr) \tt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     