A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �PNSF_SET_T   h $MODE  $IN_SIZE  $OUT_SIZE  $ADDRESS  $BY_PWFAIL  $BY_PLCCON  $BY_PLCRUN  $BY_T1ONLY  ��$$CLASS  ������   U    U�$PNSF_SET  ������U�           L    