��   �P�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�RYRUN_T   � $'�ENB 4 NU�M_PORTA �ESU@$ST�ATE P TC�OL_��PMPM�CmGRP_MA�SKZE� OTI�ONNLOG_IgNFONiAVc�FLTR_EMP�TYd $PRO�D__ L �ESTOP_DSBLA�POW_RECO�VAOPR�SA�W_� G %�$INIT	RE�SUME_TYP�EN�&J_ � 4 $($FST_IDX��P_ICI �MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI� DxMKR�-  $L{INc   �o_SIZc�x�� k. , $USE_FL�4 ��&i*SIAMA�Q#QB6'oSCAN�AXS+�INS*I��_COUNrRO��_!_TMR_VA�g�h>�i ) �'` ��R��!n�+WAR�$}iH�!{#NPCH���$$CLAS�S  ���401��5��5�6/ �055������c����\1l5�1071p5��%VA�G���<�0TP��?��A5I2.L;c ��"��	AU$��Y4d��Y34	A[2)Y3�Y4-D� &H��&GH\0pAhF	~ChF�CRhFÞChF�n@�fH�̾ChF�n@�fH��n@�&GAA4B�D!Bz08�H`0Q�Fhz0�i�Hl.S�Fyz0���H�z0��H�z0�j�H�z0�&G~SxV~P�HU@�QxVVa@2vX9~P;vXUA~PPvXa~PxvX���SxV�~P�vX��cxV�~P�vX�@%�vX�>cxV�~P�@RxV�^c(E\0P,hf=@+fhC�chf�H# �5maL�chfQ�# qfhAP{fh�D�chf�# QPhf��c�hfaPqPhf�@�2fh�# Eh�>s(Ea�@PqHvP3Fx�7nsHv�0�qHv�P%sFxw�sHv��sHvf!`�Fx1p�&G��@�q�v �s�v1��p�P�vV�p�P�vvR�p���=AD��G&�aM���U=AAP z&��^�)�����&���~�)��q�&����
&����&�ae=A����eU=A�A�&��X��@(� ��@P����P ���J.�����P@����PP���`H U��en���u ��U��U������ �F&�
n@�P(���DB���z0��?���`�����6W?05�V1 �FOLGE���U�Ue�MAKR�O'�SUCyH�eh�BIN����x�o { 2�L; 4%|�S�P��د���J{��Ʀ�U
��ǥeu$>��}1Ʀ4G�J� \�;2����`�6���� \�uu��ǥUB�� ����L?��������PA ��%�Xn@��01\0s2t_q* ����� ��!��$��&t��#tK���&�8� J�\�n߀ߒߤ�����p6}1������t)� \ttq�ttt}1�'�9�K�]� o�������%�쪣!2t� ������dss_
Wq	�Y��[�]�_tr
 ��8�J�\�n� ����������������=&��dsu	�UY[]_'� >Pbt����P����5$��� �-?Qcu��@������<����/G/Y/k/}/ �/�/�/�/�/�/�/�<���)/G?Y?k? }?�?�?�?�?�?�?�?TO��!���\2? PObOtO�O�O�O�O�O �O�O___C_U_ g_y_�_�_�_�_�_�_ �_	oo._GoYoko }o�o�o�o�o�o�o�o *oCUgy� ������	���-�8w��
d� +� -OOj�|����� ��ď֏�����0�j�� AT�BY�s���������͟�ߟ���'�9�
��N�A`�y��� ������ӯ���	��x-�?�J� ds��#��%��)j����� ��¿Կ���
��.�T@�R���V�?T�@{��ϝϯ������π��	��-�?�Q�L�N�?d�yϒߤ߶��� �������"�4�F�X�*c�V�=T�>�ߛ� �����������+�P=�O�a�L�N�=d� �������������@ 2DVhs�V�;]�<������ �);M_q
L�N�;d���� ���//0/B/T/�f/x/�V�9]�: ��/�/�/�/??'?@9?K?]?o?�?�N�9d��/�?�?�?�?
O O.O@OROdOvO�O�?N�)]�/�?�O�O �O __$_6_H_Z_l_�~_�_C�f� l�& �O�_�_�_oo,o>o@Poboto�o�o�_f�q��_�o�o�o" 4FXj|���oUf�(l�*l�,�o ����/�A�S�e��w�������`��tf�'v�l�+��� �%�7�I�[�m���� ������������� +�=�O�a�s������� ��]�Ο�����/� A�S�e�w��������� ʯ�����+�=�O� a�sυϗϩϻ���ط�P�B��t
ޏ�!�3�E� W�i�{ߍߟ߱�����ڸz�AC��D��E��F���0� B�T�f�x�������｝�t �������E��%�7�I�[� m�������������諭t!��G�H��M��N�.@Rdv �������Oǃ�"��G��Ht��M �5GYk}���������t#���I��J��Q��R %>/P/b/t/�/�/�/@�/�/�/�/�ǃ$��I�JQ�,/E? W?i?{?�?�?�?�?�?P�?�??�t%��K��L�GOYOkO}O�O �O�O�O�O�O�O_��&��K�L��P_ b_t_�_�_�_�_�_�_P�_oo��'��O�P*?Soeowo�o�o�o��o�o�o�o�(
&BO��P"/[m ��������T!��)��S�T��UM�Un��������� ȏڏ����"�o'SU*&BS��TX�U��V]�v���������П������*�5�'S+ ��Gom��������ǯ ٯ����!�3�.���,&BNt��������� ο����(�:�E�>'S-ds2 j�{� �ϟϱ����������P�/�A�L�	��.f� ߑߣߵ���������@�!�3�E�W�b�/n� ������������@�)�;�M�_�b�0v� ��������������@1CUgb�1~� ������@'9K]ob�2� ������//@//A/S/e/w/b�3� �/�/�/�/�/??%?@7?I?[?m??b�4�/ �?�?�?�?�?	OO-O@?OQOcOuO�Ob�5�? �O�O�O�O�O_#_5_@G_Y_k_}_�_b�6�O �_�_�_�_oo+o=o@Ooaoso�o�ob�7�_ �o�o�o�o!3E@Wi{��b�8�o �����)�;�M�@_�q��������x9� ׏�����1�C�U�@g�y��������x:Ə ߟ���'�9�K�]�@o����������x;Ο �����/�A�S�e�@w����������x<֯ ���%�7�I�[�m�@ϑϣϵ��ϲx=޿ ��	��-�?�Q�c�u�@�ߙ߽߫��߲x>�� ���#�5�G�Y�k�}�@��������x?�� ��+�=�O�a�s���@�����������x@�� !3EWi{�@������xA�� );M_q��@������xB /1/C/U/g/y/�/�/@�/�/�/�/�/�xC/ '?9?K?]?o?�?�?�?@�?�?�?�?�?�xD? /OAOSOeOwO�O�O�O �O�O�O�O_�u_3_ E_W_i_{_�_�_�_�_ �_�_�_o�u_7oIo [omoo�o�o�o�o�o �o�oo3EWi {������� ��(A�S�e�w��� ������я����� +�6�O�a�s������� ��͟ߟ���'�2� K�]�o���������ɯ ۯ����#�5�@�Y� k�}�������ſ׿� ����1�C�N�g�y� �ϝϯ���������	� �-�?�J�c�u߇ߙ� �߽���������)� ;�M�X�q����� ��������%�7�I� [�f������������ ����!3EWb� {������� /ASep� ������// +/=/O/a/s/~�/�/ �/�/�/�/??'?9? K?]?o?z/�?�?�?�? �?�?�?O#O5OGOYO kO}O�?�O�O�O�O�O �O__1_C_U_g_y_ �_�O�_�_�_�_�_	o o-o?oQocouo�o�_ �o�o�o�o�o) ;M_q���o� �����%�7�I� [�m�������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ư߿���'�9� K�]�oρϓϥϷ�¿ �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u�������������* _�ds
�qu����q����q�ss����tr� t�� q �t��CUg�y�������@Z��`��J L �K Mquq�s)Ars�kq) ��t!'�tt 1K]o���������A��ads����,�r8tRB,  u(H""mI Z  \9 J/\/n/�/�/�/�/�/�/�/��9��?)?;? M?_?q?�?�?�?�?�? �?�?��O%O7OIO[O mOO�O�O�O�O�O�O �OO!_3_E_W_i_{_ �_�_�_�_�_�_�_o _/oAoSoeowo�o�o �o�o�o�o�oo+ =Oas���� ����� 9�K� ]�o���������ɏۏ ����#�.�G�Y�k� }�������şן��� ��*�C�U�g�y��� ������ӯ���	�� -�8�Q�c�u������� ��Ͽ����)�;� F�_�qσϕϧϹ��� ������%�7�B�[� m�ߑߣߵ������� ���!�3�E�P�i�{� ������������� �/�A�S�^�w����� ����������+ =OZ�s���� ���'9K ]h������ ��/#/5/G/Y/k/ v�/�/�/�/�/�/�/ ??1?C?U?g?r/�? �?�?�?�?�?�?	OO -O?OQOcOuO�?�O�O �O�O�O�O__)_;_ M___q_�_�O�_�_�_ �_�_oo%o7oIo[o moo�_�o�o�o�o�o �o!3EWi{ ��o������ �/�A�S�e�w����� ���я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }���������׿��� ��1�C�U�g�yϋ� �ϯϺ�������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ �������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/�/�??'?9?K? ]?o?�?�?�?�?�?�? �?�/O#O5OGOYOkO }O�O�O�O�O�O�O�O O_1_C_U_g_y_�_ �_�_�_�_�_�__o -o?oQocouo�o�o�o �o�o�o�oo); M_q����� ����7�I�[� m��������Ǐُ� ����3�E�W�i�{� ������ß՟���� �(�A�S�e�w����� ����ѯ�����+� 6�O�a�s��������� Ϳ߿���'�2�K� ]�oρϓϥϷ����� �����#�5�@�Y�k� }ߏߡ߳��������� ��1�C�N�g�y�� �����������	�� -�?�J�c�u������� ��������); MX�q����� ��%7I[ f������ �/!/3/E/W/b{/ �/�/�/�/�/�/�/? ?/?A?S?e?p/�?�? �?�?�?�?�?OO+O =OOOaOsO~?�O�O�O �O�O�O__'_9_K_ ]_o_zO�_�_�_�_�_ �_�_o#o5oGoYoko }o�_�o�o�o�o�o�o 1CUgy� �o�����	�� -�?�Q�c�u������ ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �ϸ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy� �������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/ �/�??%?7?I?[? m??�?�?�?�?�?�? �/O!O3OEOWOiO{O �O�O�O�O�O�O�?_ _/_A_S_e_w_�_�_ �_�_�_�_�_ _o+o =oOoaoso�o�o�o�o �o�o�oo'9K ]o������ ��
#�5�G�Y�k� }�������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� &�?�Q�c�u������� ��ϯ����"�;� M�_�q���������˿ ݿ���%�0�I�[� m�ϑϣϵ������� ���!�3�>�W�i�{� �ߟ߱���������� �/�:�S�e�w��� �����������+� =�H�a�s��������� ������'9K V�o������ ��#5GRk }������� //1/C/U/`y/�/ �/�/�/�/�/�/	?? -???Q?c?n/�?�?�? �?�?�?�?OO)O;O MO_Oj?�O�O�O�O�O �O�O__%_7_I_[_ m_xO�_�_�_�_�_�_ �_o!o3oEoWoio{o �_�o�o�o�o�o�o /ASew�o� �������+� =�O�a�s�������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߲��� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASew�� ������+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ ��/?#?5?G?Y?k? }?�?�?�?�?�?�/�? OO1OCOUOgOyO�O �O�O�O�O�O�?	__ -_?_Q_c_u_�_�_�_ �_�_�_�_�Oo)o;o Mo_oqo�o�o�o�o�o �o�o�_%7I[ m������ �!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s��������� ͯ߯��� �9�K� ]�o���������ɿۿ ����#�.�G�Y�k� }Ϗϡϳ��������� ��1�