��   2W�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���C�ELL_GRP_�T   � �$'FRAME �$MOUN�T_LOCCCF�_METHOD � $CPY_SRC_IDX_�PLATFRM_�OFSCtDIM~_ $BASE{ �FSETC��A�UX_ORDER�   �X�YZ_MAP �� �LEN�GTH�TTCH�_GP_M~ a AUTORAIL_���$$CLA�SS  ��i���D��D�8LOOR ���D8�?���O��/, � 1 F �H8=_`_��D'�82 �����K!/3/E//i/{/�-_ �/�/�/pO,��p 8!�/ �/?/g?y?�?]?�? �?�?�/�?�?�?�/C?E?�13OEOWOY?�O �O�O�O�O	__	O3_@E__1O�O�O�A{_ �_�_�O�_	oo�_?o�QocoQ_{o�ogo�$�MNU>A�R�_d  8K>}��5�?�d����e�aBy�� �qC��� M�_=?Qs ������	�� �?�)�K�u�_����� �����ˏݏ��� 5�7�I�k������˟ ��ן���7�!�C� m�W�y�������ٯïկ����b!�K�2� G�i�k�}���ɿ��տ ����5��A�k�U� wϡϋϭ�������� ��	�C�-�?�a�c�u� ���߫��������-� �9�c�M�o���� ���������;�%�7�Y�[�A�1q����� ��������-9 cMo����� ��;%Gq [m������ �%//1/[/E/g/�/ {/�/�/�/�/�/�/	? 3????i?S?e?�?�?�?�?�?��A�?O�? O1O3OEOgO�O{O�O �O�O�O�O�O	_3__ ?_i_S_u_�_�_�_�_ �_�_o�_o)o+o=o _o�oso�o�o�o�o�o �o+7aKm ����������!�#�  �$M�NUFRAMEN_UM  W�>X��D  �k�TOOL A���������\ @��;��.L�K��L�����3���Ł'	��ß�	�Ær�DsF�ł��.W����K���(ڀ��ŁD�� C3  C��W���-���K�c� M�_�����������˟ 5���#�%�7�韃� m�������ů�ٯ�� %��1�[�E�W���{� ������ÿ����� E�/�Q�{�eχϱϛ� ����������)�S� =�O߉�s߅ߧߩ߻� ������=�'�I�s� ]��������겁 p�����n�2�4�F�h� ��|������������� 
4@jTv� ������� *,>`�t�� ����/,//8/ b/L/n/�/�/�/�/�/ �/�/�/ ?"?$?6?X? �?l?�?�?�?�?�?�? �?$OO0OZODOfO�O zO�O�O�O�O�O�O�O__
�13_q_X_m_ �_�_�_�_�_�_�_%o o1o[oEogo�o{o�o �o�o�o�o�o	3 /iSe���� �����)�S�=� _���s�������ˏ�� ߏ�+��'�a�K�]� �������ߟɟ�� ��!�K�5�W���k��� ����ï�ׯ��#����Y�C�U�w�y��A ��Ϳ��ɿ����!� K�5�Wρ�kύϷϡ� ��������#��/�Y� C�eߏ�yߋ��߯��� �������C�-�O�y� c����������� ��'�Q�;�]���q� �������������� ;%Gq[}�� �����I 3Ui{������  �$MN�UTOOLNUM�  
 
 �D   @!