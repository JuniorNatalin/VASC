A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DMR_GRP_T  � $MASTER_DONE  $OT_MINUS   	$OT_PLUS   	$MASTER_COUN   	$REF_DONE  $REF_POS   	$REF_COUNT   	$BCKLSH_SIGN   	$EACHMST_DON   	$SPC_COUNT   	$SPC_MOVE   	$ADAPT_INER   	$ADAPT_FRIC   	$ADAPT_COL_P   	$ADAPT_COL_M   	$ADAPT_GRAV   	$SPC_ST_HIST   	$DSP_ST_HIST   	$SHIFT_ERROR  $SPC_CNT_HIS   	$MCH_PLS_HIS   	$ARM_PARAM   d$MASTER_ANG  $DSP_ST_HIS2   	$CLDET_CNT   	$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$GRAV_MAST  E!�FMS_GRP_T t *$REM_LIFE   	$NT_LIFE   	$T_LIFE   	$CLDET_ANG   	$CLDET_DSTB   	$NT_LIFE_0   	$T_LIFE_TEMP   	$REM_LIFE_0   	$GRP_CL_TIME  $PCCOMER_CNT   	$FB_COMP_CNT   	$CMAL_DETECT   	$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $DTY_STR_T  $DTY_END_T  $CLDET_CNT   	$CLACT1   $CLACT2   $CLACT3   $CLACT4   $CLACT5   $CLACT6   $CL_OVR   $CLOMEGA1   $CLOMEGA2   $CLOMEGA3   $CLOMEGA4   $CLOMEGA5   $CLOMEGA6   $CL_FRMZ   $CLDEPT_IDX   $CLCURLINE   $CLDEST1   $CLDEST2   $CLDEST3   $CLDEST4   $CLDEST5   $CLDEST6   $CLNAME ?( �PLCL_GRP_T  � 	$CALIB_STAT  $TRQ_MGN   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	��VCAX_REFA_T  @ $REF_FACTORY  $NUM_SET  $MAST_TO_REF  $PRE_MST2REF  5<�VCAX_REFD_T  , $COMMENT $REF_UPDATE  $REF_AXIS 2 	��VCAX_REFS_T  8 $STEP_MS_ENB  $NUM_SET  $STEP_DATA  $PRE_STEP  �VCAX_REFM_T   $IS_SET  $MASTER_COUN  �VCAX_REFG_T  0 $REF_DATA 2 
$REF_STEP 2 	$PRE_MASTER 2 	�$$CLASS  ������       �$DMR_GRP 1 ������      	                                      	                                      	 ��i0� ���,5��L�3�]                 	                                      	                                      	                                     	                                	 ���� S � �S�`��^k�(A             	                                      	                    	                    	                    	                    	 ����n�����       	                   	 B B B                        	 ���������K�_�����.��             	 ��k[��������,��-�3�:             d                                                                                 =L��                                    ?�                              @�                                                                                                                                                                                                                                                           	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 �����$FMS_GRP 1������  	 G���G�H�["L0o�Im��H�)�             	 O`�,PWv�O
H�L!KHDoK9��             	 B�  B�  B�  B�  B�  B�               	 C!T�BjJa�Η�>�_¦.@B�l             	                                      	 O�pP��XO�� IQ_Kӭ�K���             	 B��B��B��B��B��B��             	 G���GϹH�^HL0o�Im�H�,�            Wl\� 	                                     	                                      	                                                                Wl\�Wl\�Wl\�Wl\�Wl\�Wl\�Wl\�Wl\�MVAcM]NXM���NFm�NFn2NFnqNFnvNFn�N�]�U%9EWl\�Wl\�X�2pX�2� 	    "                                ������������������������6��A� AϦ6�h6�6��6�6�x5�}A�������  �5$�5d�5��5��6m�6��6��6��k1���(��8�sr�x�Ȭ�ȓ��m�<9�5�  4�4�A4�e4�/4�`4�L4�>4�8 � �� �8� ��� �d� ��4 �� ��z0� �4&4�4��  ��������������������������t�����s��������������������|������  ���������������������������������0���(��(�
�7��8���;��;s�;wK��}��'����������  �"&�" �"�""�" �" �" �" ��� ȕ� șH �� �
 �	� � ���o�t ȕ��"�"%     P   P   P   P   P   P   P   P   d   d   d   d   d   -   -   -   d   d   P   P  ����������������   ���������������n��������������������       ���t������������                             ���!   ����������������      ���-��������                       ����          �����      �   �   *   ����  v����   ����  ��������           ��������      ��������      ����              ����                  ����������������    ���7�������^�������T���@����     �      ����            ����    ����       ����          �  r��������      �    ��������     d   d   d   d   d   d   d   d   �   �   �   �   �   �   �   �   d   �   d   d                                	8                                                     
   
   
   
   
   
   
   
                                    
  @44�@44�@44�@44�@44�@44�@44�@44�������bS��bJ�������k���Ϳ��f�������`��e�@44�@44�  ?��?��?��?�� ?��?��?��?��>��?��?�:>�K�>�+K>��`>��>��t?�U?��?��?��  ���{���(������
���"���
�������DZK�7^/�7`�K'S�K��K��Kk~�J1u�����6B��ā���{  ;W};W};W};W};W};W};W};W}�#�:��K:�N!�"	9�"	��!�ü!s���ck�:��2;W};W}  ���񿹟������������󿹟����������M��Z5#�Z3�F���G/�F&6�F�P�G9���9��[Y���󿹟�  ?�.z?�.z?�.z?�.z?�.z?�.z?�.z?�.z@���@���@���@���@���@���@��@���@p�@��Z?�.{?�.{  ,($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP027...........................0008      ($UP002                                     ($UP003                                     ($UP003                                     ($UP002                                     ($UP002                                     ($UP002                                     ($UP002                                     ($UP002                                     ($UP001                                     ($UP003                                     ($MAKRO004                                  ($UP027...........................0008       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      �$PLCL_GRP 1������� D    	 ?�  ?�  ?�  ?�  ?d��?zY}?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$VCAX_REF_GR 2������ t 
 �REFERENCE 1        	                                                                                                                                                 REFERENCE 2        	                                                                                                                                                 REFERENCE 3        	                                                                                                                                                 REFERENCE 4        	                                                                                                                                                 REFERENCE 5        	                                                                                                                                                 REFERENCE 6        	                                                                                                                                                 REFERENCE 7        	                                                                                                                                                 REFERENCE 8        	                                                                                                                                                 REFERENCE 9        	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE2_1       	                                                                                                                                                 REFERENCE2_2       	                                                                                                                                                 REFERENCE2_3       	                                                                                                                                                 REFERENCE2_4       	                                                                                                                                                 REFERENCE2_5       	                                                                                                                                                 REFERENCE2_6       	                                                                                                                                                 REFERENCE2_7       	                                                                                                                                                 REFERENCE2_8       	                                                                                                                                                 REFERENCE2_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE3_1       	                                                                                                                                                 REFERENCE3_2       	                                                                                                                                                 REFERENCE3_3       	                                                                                                                                                 REFERENCE3_4       	                                                                                                                                                 REFERENCE3_5       	                                                                                                                                                 REFERENCE3_6       	                                                                                                                                                 REFERENCE3_7       	                                                                                                                                                 REFERENCE3_8       	                                                                                                                                                 REFERENCE3_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE4_1       	                                                                                                                                                 REFERENCE4_2       	                                                                                                                                                 REFERENCE4_3       	                                                                                                                                                 REFERENCE4_4       	                                                                                                                                                 REFERENCE4_5       	                                                                                                                                                 REFERENCE4_6       	                                                                                                                                                 REFERENCE4_7       	                                                                                                                                                 REFERENCE4_8       	                                                                                                                                                 REFERENCE4_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                         