��  	��A��*SYST�EM*��V8.2�306 4/2�
 014 A�5  ����A�AVM_WRK_�T  � �$EXPOSUR�E  $CAMCLBDAT@ �$PS_TR�GVT��$X� aHZgDIUSfWgPgRg�LENS_CEN�T_X�YgyO�Rf   $C�MP_GC_�U�TNUMAPRE_MAST_C�� 	�GRV_}M{$NEW���	STAT_R�UNARES_E=R�VTCP6� %aTC32:dXSM�&&�#�END!ORGBK!SM��3!�UPD��ABS�; � P/   $PARA� �   ���ALRM_REC�OV�  � A�LM"ENB���&ON&! MDG�/ 0 $DEBUG1AI"d�R$3AO� TYPsE �9!_IF�� D $ENwABL@$L�T P d�#U�%Kx!;MA�$LI"��
 0�APC�OUPLED�� $!PP_PR�OCES0s!�(1Ns! h�!> Q�� � $SO{FT�T_ID�"�TOTAL_EQfs $0'0NO*2�U SPI_IND�E]?5X�"SCREEN_NAMr {�"SIGNe0��/�+!0PK_F�I� 	$TH{KY�7PANE24� � DUMMYE1d�4d!�54�1� �ARG�R�� � $T{IT�!$I�� N DdDd D�0DU5�66�67�68�69�70�7G�1EG��1E0G1:G1DG1�NG1XG2cB4�ASBN_CF>"� 8F CNV_�J� ; �"L A_C�MNT�$FL�AGS]�CHE�C�8 � ELLS�ETUP 	 �P� HOME_I�Oz0� %5SMA�CROARREPRJX{0D+>0�dR{�lT��AUTOB�ACKU�
� �)DEVIC&�3TIc0�� 0�#��PBS$IN�TERVALO#I?SP_UNI��P�_DO�V7�YFR3_F\0AINz1���1�S�C_WAx�T�Q-jOFF_� �N�DELZhLO�G�R�1ea�R?�Qf`�3?�� {1�5��<�MO� ZcE' D [MZc����aREV�BI�L�g`�AXI�� �bR  �� OD7P�a�$NO�@M�!� �ar�"w@� u<q�bZ0D�C� d E R�D_E�`Ts $�FSSBn&$CH�KBD_SE�UA�G G�0 $SLOT_�V2�q�� Vzd�%4�މQ_EDIm  _ � cQG��CPS:`a4%$EyP1T1$OP^0r2dap_OKnr;US�!P_C� �q��T�vU UPLACI�4!TQ?��p( �QC�OMM� e0$D�;�Q�J0f`�y�?�2o8�BL%0OU�r ,K�QQ2QU �B�@y O]Å���CFWt X �$GR� ��M=BZ`NFLI���0UIRE��$g"~� SWITCH���AX_N)PSs"C�F_�G� �� 
$WARNM`"`#!�!�p�@LI��f�NST� CORz-�RFLTR`�/TRAT;PTb�� $ACC�Q��N |��r$ORI��o"�RTlP_SF~g�CHGz0I��bT�1�UIʐT��K�>� x i#
Q\nr�HDR�2J; �3I�2D�3D� F�U5D�6D�7D�8D��9�"�O�D <�F �����#�܀O�_M�� t� 	PEq0�1NG�1iBA� Q���q ��!�Qp�0=q�0�I�P�PJ���F�S��pm �RC ������"J��_R��gCb��J����ļJVep�%C�X���p0��P�OF� 0  @F RO��&9�6��IT3c9�NOM_�yV�lS��P�D �0��A�B�'&�EX��B0��P��<���
$TF�E06��D3N�TO�S3�U8P+� -0PS_H�j 1�E{� %�Y#&�d%(��1}#�DBGDE}!�_p$��PU8��1a2)��I"ƻ�AX�Ae$]eTA�I�SBUFivd|Y�/ � k׶f�PI�$��P���M��M��^���F���SIMQ� ��$KEE:�PAT@0�����N#��Y"�$��L64FIX/���⥟TC_��� ����c��CI됎�PsCHOP��ADD�� �������I"m0p�3�_��!f���n!�
��a��W���d"�6$�MC�� �0yJBE�ͤz��l�+�pi���N��� ��p�CH� EMP�#$G�����p_�lS��1_FPm��@��SPE��lPn�������� V�q<r�A̛�JR�<rSE�GFRA��3 �R>�0T_LIN{sMPVFs!�$�'�_�"�#m�"� R���$�y� D ) ���`�����2�f��)P���Ţq�f�SCIZc��T����3�RSINF��G�R �e3 e��> L�з�ΚCRC(�AcCC n��3 ���*���1Ma�������D&�e#
)C+e`T�AM ^�&�T(E�VT&i�Fj!_F��N�&�@f�`�((�������'��rj1���A! �>p���-�RGB�ª�F�B ׂ��De�R��LEWر�Q�����/�. g�RWt"� ��Ư�5b��#�R� HANC�$LG~��!�QU�y�gp��6�A:`� a�c�R?2 �3p0��3�\��8RAnS�3AZ���7HP ��O�FCTC�Y07�F)����\R�ADI�KO�H @�@�o��D~�.���6�S�p����qM�PW*���M�4A�ES��l#�,�0I}_�4#  �=I+$�CSX��H�B��$*�?p�s��T�B��C�0N�p�IMG_HEIGHmq�rSWIDK��VTt��M��pF_A 8{��B`EXP�A4�N�U�CU7�]�U%�w% $_�TIT���r�s�p��E�:RZ_% {�&*�b{� ��A~�NOwPAD	q?W�i?�,�����DBPXW�O�&�'��$SqK���rt�DBT�0wTRL%�( �,��A!���@��rDJ���LAY_CAL`�q	��`�@�gPL	�~G�SERVEDW�wb�w��'��	�
��9��0���aAA%��)�b��PR� �
�`"���%�* l_���$�$"ʆ`Loy+|"�t���&�,�"�|�P�C%�-��cPENE���!.��e֠\}��r/H�0C��� *$L2�+$os��+@C�T ���O�0_D�A��RO�����䤍�|�R�IGGE�PA�US��VETUR�N���MR_�T�U>��a�EWM<F��GNAL�����$LA-��n�,{$P��-$P\@F!�.�b��C!�!��DO` ��\�H���b�GO_AWA�Y8�MOD�0�Bv�`CSrpEVIm�� 0 P $fіRB�
�PI����SPO��I_B�YT2����TXw�L$�1 H� 7��Ф��TOFB��FE�l������w�CU2��DO����0MC���N���7�`����Hry@W����  �w�wELEGR3 T����cCINKh�����5U�L��HA���}$��}  q�w�����4 ��`�MDL�� 23���(�O��^����C�2����J]�}O� m�}2�U�r�h�����2��	����
<w�%U?5� $]��0 �PcC�PZ��Pa5бw�b�ϲ��̵IDJ��˶�b˶W ���NTV��вVE��(Р$W�D�2W��J�&��<�pSAFE)����_SV�BEXCL�U�a��>2ONL���Y6��3x@�Qw��I_V�@�PPL�Y_���� Ƕ��_�M�"��VRFYI_�c��MS3�PO���x@!֧@1~S4�^�O࢐�İ��@� 6���`TA_ ����� �bW�SG�  �7 ��CUR�π�}S��tpUQO�R�EV�ٯҦ�jPUN��p��ԥ��Ё��� ��0���ѧ@���b�EFаI�r8 @b� F���T�OT� ��At<�At'qAt^�Lr�EM��NI�r9 �L �`��A�ʱ��DAY	�LOCAD��6tv�Bs5Js�EF�P$�X�:�d' SO����0��`�_RTRQX�; �D�!O��RQ{ ������:| C7 ��A;`���< 0�Z��p�Z�L>��6DU5��b;CA�� =9�[`�NSk���ID� P�W93U����V��V�_U��< �D�IAGr�u>8O *$V��T%@ep
p}R�rt��{V2`��SWB��u���R �2�;�� �OH�r�3PP2a}IR�Q}B���m������	��BA����D@�H�����=��CY ގRQDW�MS�� AZ`w0{LIFE�`�/Hq��NB�K��@��!�����C�@f�NrЀY0�QFLA�4��OV�@W.`���SUPPO�`�Aĝ��`_���z_XP�C�a��Z�W���A��B ��CT�%U? `��CACHE�'C"ۣ�կ����� SUFFI��ϰ�`%a6t��Bs6�>q -!MSW%U@� 8��KEYIMAG��TMF�C�!�с�&INPU}R w4�G�VIEL �1A �BGL�/đ��?� 	 �npfPcBMP�!g�1IN^�Tb��	UBFv�JB���d��O#Q	T�3��S��Uu59d^�;��OF��H���C �Va!gOT�F��ץ1�D[�P_GAI�Q���@�@̒��NI_�0C���5����6�PTIC��O �PE���"��}1�A{��PCF�@INy��P[E�Aq�@!� l��A$P�3D  TP��6D�7I�8T�r=�Rv�=�AVE�F�FBP�c�C���3AW_�@<���E���v�DO<4SLO��>�1TERCE/���bDL/`�J3UFU' RQ�E�e{0�P�E}1�D
�`B�FE��3N��3 qPQ;`�5�R�6�R�5
�`G�FF� 䠣�$8�Q1��G �1�0���1F����0�3�0� ��AbB��cCA#RRg#i0�9T$ <2%cyftqRD_4�06F�SN�p��T� �FSMY��DI"e�C�$�A�D��dEG�R��F 	cu0��H b�C9�0ǰY���1��@3�G dA I� { _��3]6�0 �s�1�s�1�r}� Ц$�J�z�STp@!�r)��tk��t���t<���pEMAI����/1�`SB�@AUL��K�")8}1COU�dP��}�T!���L�,�@�M�SU��IATh�RZ�U'}�N��NF SUBRT��C�p���*rw�SAV~�@� ES��m�����r��P��M�ORDM��p_RPd���ډOTT���A��P�60���s��AX��,��X�RPeYN_�>�M�b��6�௕�G3,��@IF� ����|�a=�N� �0x5��r�C_ROᐃIK�"���Ҟ��@Rp�!���8��DSP�&��PA��I(v���ä����U���D��M��pIP0Á��D } ڔTHRES�`d˕��TZۓHS�b ۓR`�E[@��V���`�@�㑤P��NV��AG����]�ؖRPFB�d���@(��!SC�bRu��M-P��FBgCMP�À�ET�aڸ�O�"FU�DU�'��QPPEP���CaDљ[���-3t�� �NOAUTO��P��$z���z���PUSy�CR���C�B�E|�w����QH��в��r�г�� �@N����S��k������������!��7��8B��9��B���1�U1�1*�17�1D�U1Q�1^�1k�2yʩ2��2�2*�2�7�2D�2Q�2^�2*k�3y�3�3��U3*�37�3D�3Qʕ3^�3k�4y�ɴO�UT� ��R � �"@	WvPRuPLC�WAR+v�`����R|�$FACm��SE��$PARM1��2m�"k���`x³�pA� �XT��N�!S <�)9I�g��0Rv��枵- F�DRdTT @ ����E-�BE8�11(OVM�4T��A\�TROV\�DT��|�MX��vP&8�{���IND��:!
���`E�PG3����� b1�`DR�I�@c�GEAR��1IOQ�KL��N�@:EFF\�k�� |�MZ_MCM1�nE4�F�UR5��U ,��V�? �0@?� Ð0��Ei@� ��p��2� V�RTP~�$VARI�5� ܻ��UP2_� W *�?�TDI�iA>�TV�� w  ��BACG��X T�p@�U�=0�)$PROGC%�?����b�IFI��� wYPa��! ���FMR2�Y ,�k��B-� Mp�1�8J\s�}0�p�L�_���AC@I�T_[U�C_LM���(DGCLFl����DYt(LD���5������P��u�Z� ) T�sFS؀�t[ P�P��":2�$EX_�!�(�!1'�נ���!53;56�G����\ ���2��4l�O�N����1�T�1Q�G�R��U��BKUv�O1�� ��PO��9�0$�W5�0�M6`LOO��1S�Mw`E�� �����`_E ] Y��%��,PM�5�^�5l��OR�Ip�1_�7 �S�M_M	�0`!IT�A/Ia�53.S��UP:P b�s -��b]$�5�v@^��G{J� EL�TO�CUS�@ONFIG��A� c1a�CrD_$U+aא�$}��A�@P� OT�G��TAk�-�3SwNSTv`PAT`�<f`RPTHJ(�N��E� ��W��BART@E`�E�p���r�AR[p<RY��SHFTR��A|QCX_SHOR1��K�.F 9@$HG�Pa>!.�OVR����P�ItP;$U�� M�AYLO0�!A��`� ���Q]���]�ERV ��Q���Z���Gv`QR`��t;e��tRC���ASYMt����A#WJ�G����E�?QkibQ�U�d@A�CU�qP�YUP��Pġ�VkOR@M��?0�1 �c�r�2�6P�@�! ��q�%d �Ƚ�xLTOC�A�1i$O�Po"����2��p�H�O��Z�REbpR`أ��)�K�Reip�RU�u}x[QDe$7PWR	 IM�ubsR_Xs8TVIS/@��b|,r�B e�� $HC!�AWDDR�H�1GR(/�$��v�R3���.��f H��S��N� ��\���\��\�*Â�|N�U��HS[��MN�!g �uB�trq�[�OL�1��h���^��0AC�RO�p�AhqND_�C1�|�a�tšROSUP��!r_ÐI1�Uq"q1��6�2��<� ��<�Q�=��<�*�<�l7�6�AC��IO���D7���G��� �gh $� Pp_D��x�0�⣂PRM_+�� ��HTT�P_|�H#�i (��OBJE���t$�LES�����ְjN0���AB%_��T�3P�S�����DBGLV1�$K�RL�yHITCOiU@�1Gf�LOC�=O�TEMPt���0��zpv{pSS���G�HWe��A#�kW�}�`INCPU���pIO�e���r������*�IBGN�$l���� 'WAI�s�aP�����R���FW	 ېLO�m��s|���y�AN�A$Bo�����p��������RTN/`��CUF_DATAp�㖠����_MG�2(/ F�>�S(SE��r�N�8REC���N�b� 2�h�I� �m @� N�_h�Y8�3t���EXEwɒ�.Ф  d_�Xu�0�}n�$SCH�`�QP�R��FLG�vQ  D2�	/�o`o�����v ��OP�8��1~�TRA�B���CS���9�p�x $C�CTA���'�IGN�M"oO҈0�M~�T�����v���vN_PC�SO�QUp��ECF Ba��Q��׀��Ғ�	�\r��L�������@D�FRs������SPTx �$���SEQ_� Z3NS��H�*�ɀ��rC�q�@Xl�S L�}Pr�Q �-@o�bc���0�se:!�IwOLN4q 8��R�$SL�$INPUT_��$�p��P- ��&��SL���!rr���#����ݐF_AuS�"s:$LO $�O��Р�r+������PHYP���^� ��<8�UOR��#t `J��(�%�s�%�|���pP�s������|������ ���UJ}R�u � 9N��UJOG�G${DI,�$J7�VdJ8O	760I�A|Xj7_LABQ�HpZ �NAPHI�� QY�D� J�7J8�0_KE}Y� �K)�ML�%v  �AVއ�P�CTRUS�F�LAG:2}0�LG�$w �����~Y3LG_SIZJ���0>� =A�=FDHI<S�1J;@ =:tsC�� �A��j�@�X_R��������5`�LNCH2x����U01#��!BpU�)!(��L2#("DAUN%E�A�)�Dtd"Z GH�Er ��M�BO}OQ�yt Bd��pIT�Ø${�e�#�N�(SCR��`�D��|[2$�MARGI�D�,�X�ct2��M�	S0�L�W�$M�=$X��JGMC7MNCHL�M�FN�F6Kl7q�j9UFx8�Px8n�vx8HL�9STPx:�Vx8àx8� x8RS"�9H�`�;U�C�T�3 �bX�p7CIU䑌4@7�R,6� +�2G\9lPPO�G�:�%�3Ԇd2OCG�{8���GU%Ij5I�3�B(3 S43Sh0l1�P�rC�9��&�P�!N݁-�A�NAM�Qq�QVAI|� �CLEARfDn�HId�~Sr�~R5O�XO�WSI�W�XS�X8lҸ�i�i1���Tքn�DEV��}8�!_BUFFq�z� �pT0R$�IEM����' Q�
bjqq{� �pp���ˁIpOS1jeu2je3ja �
b~Q	p| �! ߈�a�ZS��{���IDX�tP�ƞ@z�jK�Tʤ�Re Y���a /{$EvC{T��v)v �"�!�} L�s������`�����w3��u(Kc~�#_ ~ �� +�#��!�s��M�C" �! C�LDP��vUTRQLI� wT2 �y�t�� ���p͑�nQD���ڠL���t�ORG2 B!�'���������!�p�s͔� �����tE�t�SV�_PT�p��R�Ǆ>φRCLMC݄m������MI;SC� d%!�a�RQ����DSTB��` K��!X��AXvR� [�t�EX�CESm 8R-�M��⡂ ?��vT �-��㠃
�M�_�I������r�����MK��c \�P�MBۢ�LICL�B� QU�IRE,CMO>�O�N�DEBU���G�ML���Ш���e�H�Pށ�ԇ�2�Di $�D�$U�PyACKE�D����DPxv��IN�b$q�_Q �pI� U�������/�	��=�U�4�T�I�ÐND:!SSb�#""$f��DC�6$IN]ю3'RSMD ���PN�r�BC��y�P{ST��� 4q�;��fRIl �e�e�ANG�bI�����AQ���;�$3ON,"�MFq T��i��00�uz� 3��SUP�� H��FX&�IGG�! � �ဃs��#�s6F�tR{�v��b������ȵ�����+�DAsTA���ETI8 f,�h1�1`INb�� t?�MD?�I�n!)M���YӇ�U�H8#�SX�DIA�Y�ANSWe�Y�Pa�A:X�Dl#)�1��ŀ��� ��CU�SV���I��&��LOf �������&G����5������ � d�MRR}22��� ���J!Á d$C'ALIQ��GrQD�2f`RIN�0G�<;$RR�SW0������ABCS�D_J�2SEe�I�L�_Ju3��
��1SP$m I�P����3������I���J�����āOaIM��CSKP�z<�- kS<�	Jm!�Q<�m�S�m�c��_AZ˂	���ELa���OCM1P&����1�� ��F�`1���� ��Z����INTEVpBSb���2I��Vp_N���7�a�'��3̒�A	DI|�����DH��t6 ���Y`$VQ�l���a$l1$ `�!`��Q`-��2��H �$B�E���	�qACCE�L����� IR�C_R-��ONT<�a�c$PS���rL  �!�s x-!sPPATH�	�Z�Z3)����_@ga���ʂ�C���� _MG�Q$D�D��"$FW�5�1������D}E�PPABN1ROTSPEE��ka/�pc�kaDEF�ۑ�)$USE)_P�>SP�C�@>S�Y
 � ʁ �aYN�1�Ac�x&,�o�x!M�OU�NGtB�O9LJ�$INC�� ����X��'3�Y�ENCSP��I�!�V�IN�bI)52Ќ�c�VE� H�*22�3_U>��<3LOWL�Qz@���p�%\6D]@I�3� �p�%r�C' #6MOS�P��MO���`ʇPE�RCH  y3OV p t"�7�a�3��_2��������b%��P*�A)EL=T*��)�$5p��_:ZFu6TRK�4�bAY��Cܑ�A)��E�C!��`�RTI8���"�`MOM�BX�@ܒc���G��D��C�\jb� DU2��S�_BCKLSH_C)U� �6�0�#���:T�"EZ�!e�CLA�L2`"2���@�`wUC�HK�p�eS� RT	Y���5$�U�0�9_�c�4_UM���Y9C�S�SCL�T# 7LMT��_Lg����T�gE m!`k�P e��0Q�!&@bd&�8PC�1�8H�pl�d��UC뀎rXT� .�CN__�N���f&�SF��9Vb""��7��a)u�hCAT�^SHo�_���& U�Q6��*����3PA�T�"_P�U�C_�p�P�F�0�q�C�t��UJG�����sJ0O�G�g�BTORQU T ��3�I�/��2�A��_W�E�D���7��6��6�I>�I
L�I�F9�)��,#�VC� 0R�䒂��1����Əc���J�RK�������DBOL_SM�!5BM���_DL�5BGRV�=�6��6���H_p���]d�COSq��@q�LN�������� � �� ��h�Қ����b�Z���6�MY����}�TH��1�TH�ET0e5NK23��[����CB`�C5B�CT�ASƱ��`h������`�SB����k�GTSE�#!C��� ���|s���ϓ$DU�P>G�D��!����3��AQ��&�$NEB��I��#���L$~ O�AS�|���8c�n�n�LPHq�Z�45Z�S��ͳ��ͳϕ@Z�ޖ�����~ V��QV��� ��VźVһUV�V�V��V
�V�H�����µ�:qT��һH�H�H��UH
�H�O��O���OIٴ�OźOһO��O�O��O
�O��FZ��������ԑ��SPBALANC�E�~aLEȠH_S�SP��4���4�>ϖPFULC8�_�G�_�ϕ!
1���U�TO_�P�uT1T2���2N�Quc� ��O�Aa�?�0��A�TK@O���'�IN�SEGu~1REV8B�~01DIFtEF	�1�+�r1�IPO!B!�gQ@��G2�����Q�LCHWAR�
"g"AB�q�E$MECH�� ��!���VAX�APEd��u���� 
����n5ROB�0CR)����b S�MS�K_��� P ��_R R���+:!vD1r/0-"+ ,3�ET+ �IN��MTCOM_C��>� �  �3�~ !$NORE3>��OPWO��� ߗ, k SB5U��QOP� ʿT�
U�=PR�UNq�PAR Dp�����0_OU�!��S�AB�"$^ IMAGVQ( �B�P�IM� BI�N'�BRGOVCRD<��	@P!Ap!_��q��R��`RB�`��[aM�C_EDT_� �K`Nl�M�JaPMwY19Ia�n�SL6�" � x �$OVSL��S;DI0DEX�c&H�cKA "V�!$N'! �5 %#:'5(����_� �" � @�@l"���2� �2�
&_���'�!�! w��0�ECT�  � H(��P�ATUSP{@C�D�ZDX�&BTM$�'�!I	�4Ia�#\�" � D( E�"�"Z�E4��!FI�LEJ@gP�!EXE�� �Q�72K24t#��{ ) � UPDATfZ1$T�HXNDP�������9p�P�G��UB��!���!�!�#JMP�WAI'pP*#�5L	O`�F�p�!��RCVFAIL_C�A��1R�@� �V��a�d��<E�R_P=L�#DBTB�q�U'BWD.F� U�P/E�IGI��TN1L#p0D�BRT�� �ERVE�c�D�b}h�1DEFSP�P � L( ���@p``�qp�CUNI"�7�@�1RR0!�.�_uL�P�! �0r !� 0�q�!N] ATA$�uNP�gKET$R#�BUt�PIPB!� h~�ARSIZEp�@E0GQ�RS� OR~�#FORMAT���uDCO�Q�EM2���TSUX� :" ��PLIpB~!�  $| �P_SWIp������U@p@AL__ � $�AAV�B���CVD	�$EZ1�`C_�zA� � � 1Q�VaJ3��V�80RTIA4hi5�hi6VMOMEN�Ttc�c�c�c�c| B @ADtc�f�c�f�cPU��NR�d�e�c��e�b ��S�P H$PIQ� �6�H�Z�l�~���! ڦ������ ��GQ�&_SPEED�G�R �tE�D�v�DE�,@��v��x��y�ESAM#��F��wL�EMOV_AXI�! �z��%���7�z��@)1d��2dR	 md`��	`a Б�INڌ 	`/����؄B�#�x��#�C�GAMM���A��R��GET�rF�IMS�PDcd
��L'IBR�1�BI�@bS/$HI�0_^� $f��E`ŘA���ӖLW�� ����$� Ӗ?b���@aCfEq��|�  $PGDCK����_.��PdւSiaɅ���c���f��c W�$I� R��DW�0�1"D��LEa�qЫ!�?hᠣVpMS�WFL1DM`SC%R�86�37+�U��q �S]�p7�P��URB����GR��S_SA�VE_D����3NOC`C�!�2Dd���� Sj<v幾Uy�mpʀ���pW�v<Ƚ�.aO�AA��񊅰���e �x��vv��ǜ�Z�\���1 ��QMuߦ � ��YL 5s~�ɇ��~�����N$B�����WѰ�(��4��`�����M��L�CLK�aDi�^�1j��P�M�� � � 9$���$W�Є�NG1]a��d��#d ��*d��1dV@��s��(�S��	`XPO+ca�Z&��P@t� p�| ��Uv������,�;�Ca_�� |�Si���i��c��@�c��mj	���jE@$��f!x��y��'Q^`���P�Q�PM4 Q}UP� � 88PqQ�𽡤QTH� sHO��HYS�P3ES����UEr��hP��� � @6B;Q#��#��_� 0'Ѵt���EN/	PBG_@B�[mB?�H#*#Jہ��I��pEW �vGTF�-b"�PO�4��   �𮗫"UyN� N� �{ �rp� PD�E���-3�BROGRA��!�264M ��I�Th@�{ INFO�� � ����`� (v�SLEQ�v6�u�6�p��D�0p�D����Ov����#���E��NU��AUyT���COPY��P�0��qʰM��N���^�PRU���� �gQRGADJv!�2wRX'��B$P&3�&W(P(��$��s	 �3EXF@YCn���!NS�T�� �4ALGO�k�.`NYQ_FREQ��U �w�!�T�LAhC�!��b.��5�CRE�0��l�IFlQq�NAT�%�${_GhCSTAT�@4��M@R���31	����Q31��|$ELE��0 �Nb�SEASIr1���"�a2 �1���6BƀIa�"`�q��M���2AB�Q�/`E� �pVU1�6BCAS9b�5����U�@�� ��$�1FV��|$��� X ~�2 2� 	� ���QFBPGQ|р�9eE|F dT|$P�Fe1�=GRIDd��SB|P�wTYs3;(| OTO �1Q)�m�� _4!E �B�wRO$��$� �v��LI:�PORAS��C'v�BSRV0)lTVDI�PT_�p@6PHT��RW�pRW4PYU5PY6PY7PY84Q���PFs�e1�~� $VALU�3ȕ��4���R�$��| n5	��C
1���0AN���R1�Rp�!��TOTA�LQ���7cPW�#I|�AMdREGENKj`b4�X!G�s�&��f�m�TRC�rKa_S���g``�3V'����c>�1E:3�@��ܚcV_H�@DA8}��`pS_YƱ�ڻ&Se�AR}�2��>@CONFIG_CSE��`RJ5_� ����Q�E� 4�{�O�v�k�F�PSܢ�F�f�C_YF��m���L�����(cMϰ���q�rd^⃁z��DEհ�"�KEEP_HNADD�q!��0�	CO�0+��A�r%�,�Of�
���q�,��1��,�REMC�@+����Bh����U4�e+�HPWD  �q��SBM!�p�uB� ,v�F1L�з���YN�p�M:�C���pQ�Er�� �l0DB�M�TRI�DA,�Bx� 0�K�TCLA�����U AYNSP��֡SEAꠁ�GK_P�Tn���B���RGIn�QSOL!UK ��P��)a&�$SC`0D�#ے�ALI�r���S�p�B#U�A}������� ���w1�q_�P�H�TIC�[�`�p[�REVIo��OLP���p��FK��_F�SSE�GQ���b��ITc3� �l0CP���TU� MSEC��MN���̢���H��`�0�G����0O��1�$N�̡_�e�$�PA� j�P�vO�iP��MLr P�<� ~�  ������e1��  $#OW-����G�����p���Hp2C�ĹAPü�!ߤX�AX�Q��A7HI��6� �ٔ�2��Ϛ���BV�EP���P�`Q���H�ߢ�r
��V�t��`a�B ^"$4:�Q������p��M��y�O��l""�S�MH��<�M=�2�� ��WRUP�_DLY��ÆDGELAk�>a2Yߔ��� ,�QSK=I'�� �P���O��NT\P�B��P �����`
��P���a ��v��l���vP�ڃP��ڐP�ڝP�ڪP��9N���J2#����yrEX@T�#z�����z�.@�z�����RDCa�� � ��0TORq���	��!�����SDRG��H��k���1Gg��eER�qUB�SPC�G�z�?2/TH2N�!D�#�?1� ���@��;11�� l�p2�F17��Ta��� Oѯ%��^������SD��VAHOME��� @]�2e�� k�}���������.�]�3e������0�B �]�4e���ew���� �]�5e�����*< �]�6e��_q����W �]�7e����� //$/6/�P]�8e��Y/k/}/�/�/�/��Sπf��_��A1X^�u`� V��-ET�yp��m2L.fk3IO�p�:I0Գ���R��W�� �� U0K�����(d ���2$�DSаIGNAL�#gf�CJ�1���RS232q5� Ɍ���%8��IC�Et����³��IT|q&aOPBIT"coFLOWCpTR00�3b��UXsCU+�MN�SUXTđ��I���FAC1Dų%@ ��	@CHQ� @h{p�p��C�$�`��`OM,p_���ET\ޠ�sUPD�pA3� T	@P�@�Qկ� !�(s�A������)��.�ERIOc��PT:p3T�2�_���Q/PDAMVWR���/9D��qV��6?FRIEND(�@��UFi��t�P���UM�YH�p@���GTHo_VTE�TIR����R�P�XUFI�NV_��ѥ�WOAITI���WX��l�Y7fG27WG1� �@1SQbbgpp_�RE�O_t��s�Q�`��[PqC�C�u��_TC3�8�Ķp�e��GˀŲ
tqֱ@&Q/A�r�j�QX�EV��Ea��������D�X s�ML����`��SXP��]E#T�CG3�WCP�gws�|tD�LOCKkuvӮ�V��q�t&a�$�f[���pkQ�e�qY1}XlP2o[2
�{3o[3}Z�y'�~Y��yC�6.�s.�r$)VV��V8eVl��Q��a�b!�غ��F �sρ��fqB���`�Rh�ɠ��E�$߂��S�@a�Tu���PR����uj�Sl�G��2f0�D�� ����D%s[��w���[���p��@|`�@��
J �BS޸1� ؚ�R_�6�oQ���`RUN���AXSA�`A�PLX�QV⮒THb�J�X��6�aqTF"�NT�>��IF_CHeS��`~�qU��6��G1���0���� 6�_�JF?�PR�`���{RTC� ���gGROf�A�MBVqb̐CrÃ��`UI#�v��BU)cRSM}���a`r�_W�P�ToBC_P�PCM��9D��ЖLDR��ރ��A��@��c�ITl�"�� ���TA��G� s���|� ��ę��� ���� �ݾ2�  2� ��S��g��	|# �Vд�}�I�t��ˀ~�TOT��~�D|젖�JOGLIzCN
`E_P��qBO���}����`�FK��_M#IR��Ѵ{`M>r�AP]q��E)P�Ҕ�J�SYS�˂J�PG'�BRK�bѕߐ:��I"1  N�pS�Y�x�D�A~��B�SO�}��0N��D�UMMY15U��$SVVpDE_O�PoCSFSPD_�OVRU��� L�D��óOR��� N�P��Fߑ�Ʈ�OV���SFڟ��.�F� �́ճc8ؿQ˂L�CHDLz�REC�OV��[P��W�PM��vձ�ROoC����9_ ��� @�&`�VER��$OFeS&`C;��SWD���r�����Rū�TR��1W1FpE_FD�Oƃ�Ӡ��B��BAL�����1K0%�V�A �B�@��b� �G�,�AM*Ã�D�Z��t�_M0�|B��3��T�$CA���DU����HBK�AЖ��I�OoU��1qPPA�����������2~��DVC_DB)c�0�ё�21���́H�1�P���H�3P���AT�IOˀ�A{���U8tS젆6CAB��nR��c7p���`S��A��_��@ЖSUBCPU�2��Scp�0�B��@�sj�B��2��$HW_C_ dЧs5�sAta���$UN�ITb�\ U AT�TRI�i��CY{CLϳNECA�����FLTR_2_�FI��8���6��Pxǻ��_SCT�cF_UF__�q
�FS�1:�ZCHA��Q�)9�qB(RS�D���2x�ޣ�1�0_TW�PRO����g@KEM*0_��V�T�q� z��D�IPҔRAILAiC>��bMg�LOu��S��9�R܀��䁟�V��PR2�S�a�p�!C$�$@	��FUsNC���RIN�`0Ԥ�'$fARA8 �b� ��P#X0��P#W3AR/���BL�af'$Az+v}(v(DA``�Q!�(�#z%LD�@ ��q�#��Z!ہ�#�TI�5y���$��@RIA�A�2AF
��P;A.3��45�p8�r@�MOI` �ևDF_�P7��Ac�L�M��FA�PHRDYJTORG͢��fS|� �5MULSE�P�����J��J�������FAN_A�LMLVV�AWR=N	EHARDpP�E��Y"2$SHADOWl��/�?Bc�@�w@u�:�_m�ЖAU��`�:�|@O_SBR&�E���JU &�/!��CMPINF��pk�D�!�CREGpUq��л�i�� J�v�Q$;Q$Za�e�O�j��� ��EG�~���*Q#AR�����2�q7Wܧ ,�AXE��ROAB��������R�_�]�w�SY_�dQU��VS��WWRI�P=V5 SCTR����T���EW�8�FT�qkB�`B��P���V,�����OT�O�A8���ARY���3b���B�ƱFI,5�ܳ$��Kq1��JSa]�_�S��EU:3�zbXYZ'B�j�5�fOFF��Rb�zbnh7`B��"`�d��V�  �cFI� ��gq��«�"��_aJ��6���y�$a@ddk6�qTB)qd�2arC� �DU�ҺDV7�TUR@X
3�uAa�BX�P��IwFLg�Tд�7P�p�ex�Z�û� 1�8�K��MДDV����ORQy��V#�W3I��2�+�s0��h�à�Tz�OVE����M� *��C��S ��
R��6@��*A��W  ��<�! �50����� ݀Q�*�������'�S�'���ER��Z!	B�E�PD��e�A����eH%t?g�!���!AX��6��! Ua���˙�1˙�`ʚ �`ʚZpʚ�pʚ��ʚ�ʚ1_�ʖ�0Ǚ�0 י�0癮0���0��0 ��0'��07��0G�d��X�DEBU-$�(!4C����vbAB������~�V��, 
#�Y�?�K�OW� #aW��aW��aW�ZqW� �qW���W��:4fp42\���cLAB�bI�) 6�GRO� Ir-L��B_�L��T�� �`�@ �4�J�0�A<�AND���Z���e]�Ay� ���@~a��0�!�ȡ ~`NT@=!?�SERVE��P�� $�pT Ae�!��PO��K@��-`z��0��_MRAQ_� d � T�Ўe�ERRr2�00T)Y2�I��V�`��N7�TOQ����LhP8���RJ� ���D@>Q � p��4��Ԯ�_V1f��������2��2���D@��p�H����$WT� �֘q�VQ��@�$���d0��|���OC�!P� � �COUNT��Q ��SHELL_CFGQ�� 5!pB_wBASVCRSR�SAB� ~SSWT�!h�1��%g�2��U3��4��5��6���7��8��[�ROO0�0��Y`}`NLQls�AB�úi�ACK4�IN�T� ���0pa@�0�_PU�,0@�OU�3Ps l���I����TPF?WD_KAR<ї0&�RE�Ę0PO`�! QUEr�t��� �r.@_AI@7�H�{`p�D��EzbSEM?`Ox0)6�TY*�3SO��)�DI6�s p����b1_TM��N'NRQg{`E� �(�$KEYSWITCH���I��{HEupBEAT�qE:PLE;���U��F���SND_O_HOM20O<#7REFe�PR�a��(�Q�P7�C� O�1��v�O �;rK@0IO�CMgt��a� �G�HKQ� D<xat�RESUUB���M�"��w�wsFOR�Cx�#\�G�O}M;P � @�T*3~@U�SP9P1��$9P3�4� ���S�HDDN�P� �BL�OB  �pPNP�X_ASP�� 0�v�ADD�GA$�SIZ�A$VA�:���0TIP��'#�A�� � �$c�( �`bRS���"QC7Л&FRI	FHB�S���� {NFjODBU�P����%�#�)�� �s�Si�P� x��SIT�TE�sX��s�SGL#1Tab�p&���<3íP$0STM�T�qU3P&P�VBW<��%4SHOW]5�A�SVDTU��; ��A00~Ħ2 ��7��7��7 �7U5�96�97�98�99�9A�9\P�7��7 ӱ�6�P�7�C�3W�pH��91�91�91�91��91�91I1I1� I1-I1:I1GI1�TI1aI1nI2�92 �9`@X�9�`@X�9Yp�@XI�p@X I2-I2�:I2GI2TI2aI2PnI^�h�93�93�9U3�93�93�93IU3I3 I3-I3:IU3GI3TI3aI3nIU4�94�94�94�9U4�94�94�94IU4I4 I4-I4:IU4GI4TI4aI4nIU5�95�95�95�9U5�95�95�95IU5I5 I5-I5:IU5GI5TI5aI5nIU6�y6�96�96�9U6�96�96�96IU6I6 I6-I6:IU6GI6TI6aI6nIU7�y7�97�97�9U7�97�97�97IU7I7 I7-I7:IU7'�7TI7aI7nD� @ē0P� UP�D���"+���
L��0GUN_C���� `�g�PUT�'�IN\���<AX�|�GO�U��G�I��IO_SCA�w�0YSLOP�� � E%�"#��' :'� d�� ʤ	�PԒ� �R��F��ID�_Lj+�HI&�I���LE_g�V���k$��SA���� hЂ�E_B�LCK��M1��D_CPU��F ��: �&�Y�k�Է��b�Rw ��
PW"��� 	�LA�2S������RJ�FL O5��5�đ 8�V���V���TBC�#�C!�X -$}�LEN��$L}�D�RA��d!$���W_��&�1}�C�2���M�b��� 3�I�I� ]���TOR���}��D����� LACEG��}������ _MA+ �J� ׎J�TCVQ�r� �T ssڒՈ�����d ���JF��$M��"��J���0��� ���2/ ~0����6��JK(�VK:�4$B�3,�J0O�>��JJF�JJN�AAAL>�t�F�t�n�4o�5��N1�ܥ�d��N�y�L��{� �6x�CF/!�T�v��M?1�"B�NFL�IC�# REQUwIREEBUO�y���$Tx�2��6�z� �x�. �3�{ \rAPPR,�iC��{�
��ENs��CLOS� ��S_�M� $ ���
�$���A?  �����  ����%���������s�VM_WRK� 2 ��� 0  �#5��)L L	#�`�����!�q���_� �n�+5U 1;M_��� ���/B/T/7I+ k}�5/ �/�?�/-?;?1/@r?�?g/y/�9&�D�/ �/�/e?O�/6O?O?�]OkOa?�O�O�K��B�SPOSU� 1���� < �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ����
���B~�N�L�MT�����C  �1�IN:�L�0�PRE_EXE]�1��l�.�AT}��J�����LARMRE?COV ��l���DLMDG � "�LM_IOF ��d� *�<�N�`�n������x��ǯح, 
�O����FNGTOL �!�I�@A �05�C����PP��N ?��������Handlin�gTool �� �
V8.20Pg/A2E�������88150�������
33477126��� ��Ű������葿��7DE3����	F�.014i��FRL�����2���X��TIV}�l�J��i�UTO�� ��h�P_CHGAPON=���������L�1	� @��������I��U� 1 f���>j��4����VI�Q�c߽߇������ �{����HG�����HTTHKY�ߚ߬����� 6�H�Z�l�~���� �������� �2�D� V�h�z�������
�� ����.@Rd v������ *<N`r� ��/���// &/8/J/\/n/�/�/�/ �/�/�/�/
??"?4? F?X?j?|?�?�?�?�? �?�?OOO0OBOTO fOxO�O�O�O�O�O�O ___,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $`6HZlu*�TO��uχ�DO_CLE�AN�ϧ��sNM  #��9�K�]��o����_DSPDgRYR���HI���@(����%�7� I�[�m��������ǟ$�MAXZ��t�q�q���X�t����i�PLUGG���w�î��PRC��B�"ϋޏП?�OD���^��SEGF��K�� �����'����%�87�o���LAP̏߮ �Ӌ�������ӿ����	��-�?�Q�cϨ�T�OTAL�0���U�SENU̠�� �x���r*�RG_S�TRING 1~��
�M���Se�
��_ITwEM1�  ne� �0�B�T�f�xߊߜ� ������������,��>�P�b�t�I/�O SIGNAL���Tryou�t Mode��Inp��Simu�lated�O�ut��OVE�RRɀ = 10�0�In cy�cl���Pro?g Abor������Status��	Heartb�eat�MH �FaulD�M�AlerW���u���������������� �s���q�hz �������
 .@Rdv���.WOR����� X�//0/B/T/f/ x/�/�/�/�/�/�/�/�??,?>?P?b>PO��8�0�q?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O8�O_�2DEV�>,P �?_S_e_w_�_�_�_ �_�_�_�_oo+o=o�Ooaoso�o�o�oPALTD�a��o�o 
.@Rdv� ��������8*�<��oGRI��� t��oN�������ҏ� ����,�>�P�b�t� ��������Ο��b���RD����@�R�d� v���������Я��� ��*�<�N�`�r����PREG�n��0� �������,�>�P� b�tφϘϪϼ����������(ߊ��$A�RG_�D ?	����k���  	]$��	[�]������^�SBN_�CONFIG �kۊ���CII�_SAVE  �������^�TCEL�LSETUP �j�%  OME_�IO���%MO�V_H!�4�:�RE�P���X�UTOB�ACK�
���FRA:\��� �調'`#������ ���x��15/12�/04 02:0/1:34���ت�`B�T���x��숄�����������"��� ��Pbt���5 ���(:� ^p����C��� //$/6/H/'���  ��_��_\A�TBCKCTL.�TMP DATE.D�l�/�/�/�/��INI�`��֞�?MESSAG���!���s�����1ODE�_D&���?E_Ox.P0?��PAUS�1�!�k� (q7n҈?�;)�?��?�9�?�?�0I|�?O��(OO 5O#OYOGO}OkO�O�J�c4m0TSK  �s=���/��UPDT�'0�'dP5XI�S��UNT 1|k��� � 	�@�����"���.݉bE�X-c����GQ=/ `�1� Xm� ^�&� 4�{ a�u�b^�_�_GP80� 0��zХ��=8 K�<O��8�_����_�_!ooEo0oio To�oxo�o�o�o�o�o �o/S>P� t������� +��O�:�s�^�������������\�)QME-T�15]Pޏ7� ڏ[�F��j������� ٟğ���!��E����SCRDCFG �1k�������@����� ȯگ�����"���E� W�i�{�����
�ÿ.� �����/�A�SϾ�YԤ�GR.PPQ?}��j NAN�j�	ܤ�z�_ED� 1�t�� 
 �%=-p EDT-k�b��FOLGE011���/�� @�-(����/�����?��Ϛ�  ����2���a������Q�  9۹�$�k��ڴ�g��a3\��ߩ��;R <؅���7�}���m��!4(���u������Q�@������9���5��  ���Od��������w��6�0 Tf�T��C���7��� f�@ /gy/���8X/d��/�.���/�/ 3/E/�/i/��9$?�/q?�/���M?�?�/?�?5?��CR���<O NO�O�O�?�?qO�?�}���NO_DEL��ϛ�GE_UNU�SE�ϙ�LAL_�OUT �� � gҜ�WD_AB�ORT
_{�CPIT�R_RTN  �/����CPNONS�TO��nT ����$CE_OPT;IOkX�ƣP�RIA_I	PnUԶP���PFn��+[ڳ%��Q_PARAMGP 1+[�^g�Qoco�uo4kC�  �n���`��`��`��`Ȫ�`Ҙ`ܘ`�`�`�  D�`��`�`�`�d�ؘ`�m�a	��bD"�p/�`;pH�`T�pa�`mpz�`��@ D�p�� D�`/�?��o>og�y��n|�`��`���`�� C��p���p��p��p��`���`��`��`Ř`ʪ�pмpּpܼp�
�p�`���� �|;Mv�������� ��1��ŏ׏��� I�[�m���������� -�?�Q�����	���i��PHE�@ONF�IGK_��G_PR�I 1+[  �խ�د���� �2��D�V���KPAUS?POS 1���S ,]E������ƿ ���Կ� �
�D�.� T�z�dϞψϮ���j��O�Q�_�7�QO�_MORGRP �2l ��0-A��Odr�:� 	 :�R�@�v�dߚ߈� k�������������2� ���h�V��z��:� L�������
�@�.���c�!݋���? o�o��`��0K���1r�����������������PP��+U��` UaÃ-��k}��:
 \�	�0P�N@f���5�`�53D�B��+YI�2)cpmidbg�[@m:�  !!>y�RApG��k�`�������E���`��P���-/�U��0֒0��g/�v/A/kPO�f�e/�/���/?ud�1:�/?�7"DE�F ��7)��!c!buf.t�xt?e?4 _L�64FIX , ��?�\�? �?�?�?&OOJO\O;O �O�OqO�O�O�O�O�O`�O"_4_F_~?MC�u,P  d�_P�_�UfS�t]��T|�Ub=P��Cp�Bp:�B��>B��M�B�ڢB���B��C�=!��
;�C�:��C�2RC�c�*DVP�C�H��Dw3�mE���zE#�WE@��Fu�E�?KF����	r����]��YT_�o�o �o�o�odovo�o�oO :s^�*� ��� �9���s�2:g� =<�	�%�����, 3�[��� x,��a|C*<�0<��<�p  D|mс�D��D{l��E�π�  Em�s�⁾πl)E�3� F�E���fE��fL�� � >�33 ;�I�s�n,��@s�G5�Q���� A��UL��<#�
��2����/����~`���Q���Q��E��� � H���1�9�#J;#�H�2��Z�� J�9�Q�e�w������� ��џ���B��f�=� ��a�s���������ͯ ����'�t�s�]� �ρ��ϥ���ɿۿ���5�#�v�2RSMOFST 6>쵂�9T1�PDE 3!=�pG���;�3�U�O�>/TEST02���R7"r��|�| CC4�ʀ��� ���!�Cz�P���R���sC� i�-J:�d�
-�I_1�#�7�-�T_00PR_OG %r�%v?���*�T_INUSER  ��(�C���KEY_TBL�  ��(���@0�	
��� !"#�$%&'()*+�,-./0123�456789:;�<=>?@ABC�00GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾��������͓��������������������������������������������������?������t����LCK�����S�TAT`+�_AU/TO_D� �%��INDT_ENB�� ��П�Ty2�-�STOP���SXCh� 2$�B� 
 8
S�ONY XC-5�6L輸ࡀ�@���ʹt( А;OHR5ƀK�ȼ�o�7��ACff���// � >/P/+/t/�/a/�/�/ �/�/�/�/?(??L?�^?�TRL��LE�TE� �	T_�POPU��-�T�_QUICKMEyN�4SCRE�0�B��kc�sc�4��0�9��Wc_�4UM�0�U 1��  <K�%k?gOK�EO �O�O/ÁO�O�O�DF<���_�O_P_�LS�tart SM �Comm %IBSCMANS[_�NEndxV�@�U��0�_�]User �Cancel�RU?CANCAC� o��L
�RReset>�BURES oo 3_E_�oYoko�o�o�o��o�o�@Zang=e�GZG_-A�_ �ocuL^�� �����)� ���_��ZVAG_KO�NFIG.�RVW�)��=�O�؏s�-D�ateieL�%DATEI�1��� ��E��.�@���d�v��ß������П"bMa�cro Step� tt�PMSK_�}<��LWait� Monitor3aSHTP�G�L��柫��������ZC�YCLE POW�PPWD������ DOW�%	>#�_MAINu�a�<%Cb�NUAL�?�7ZCD��&��C�[�	��������?�|(��$DBC�O� RI�Ќ5#D?BLOVRD�%ǿNUMLIM���d���DBPXWORK 1'���ϩϻ��������DBTB_1 I(7�P�Q���s�DB_AWAYý�GCP ��=��3�_ALU��?3���Y�5��$�_D�BG 1)�� �,I��,����
��
�߶�ޟ��r�%M� It�B�@��	��ONTIM�7�&���)��
)���MOTNEND����RECORD ;1/�� �����OG�O�����ٯ��y������B�XECUTING

 �~ �@	����)�P������������{E�����Q�@����/���������Ԃ������b��Pb��q���������Ϊ��͌��S����v+���#��ϝ�҂���ҏ����`��=������$���J��L>�#Kn
��  ��b��//A/S/��w/����?V��@��
 @?������/�/�/c/?�?���@���B�6���QELLED�(� )?�?�? ?�?�?���?��B���&O8O�?�?nO�? �OO�O�O�O�O�O_0O4_�O��|[��f_ x_�_�O�__�_A_��p��o)o�_Mo8o �_�o�_�o�o�o:o���TOLERENC�@�Bȉ�N�L����CSS_DEV�ICE 10�  &ƹƹWi {�������|��sLS 11,} F:E�W�i�{��������Ï�PARAM C2����TuTut�RBT 24,|�8��<I�� {C�vd ¦�s�HR�&���S�h˴��?�k۶�pm�&��\Z�g@��B˴��A��J��p�t0�pɎ��?�B�삗Ʌâvgĸ`���\�7�1����p@�Ɉc��Ɇ��� Z�l���������Ưد��7�� �m��C���Dzd0�����ѰB��A_ə�AU��������B.��Ɋ4����B� B�p���̱C"��(p�}��[33BD����ff��¿Կj���a� �G� X�( X�� Q�� vy�Ɍ)� K�]���E�sυϗϩ� �������>��'�9� K�]�o߼ߓߥ����� �������#�p�G�Y� ���3���������� *��N�9�r���_ύ� ������������8 !3�Wi�� �����4 jAS�w��� c�/�0/B/-/f/Q/ �/u/�/������/� �/�/>??'?t?K?]? o?�?�?�?�?�?�?(O �?O#O5OGOYO�O}O �O�O�O�O�O$_�/H_ 3_l_W_�_�_�_�_�_ �_�/�O_2o�Oo-o ?oQoco�o�o�o�o�o �o�o�od;M �q������ ��N�`��_��o��� ��̏������&�o /�A�n�E�W���{��� ���ß՟"����X� /�A�S���w���֯�� �������T�+�=� ����������Ͽ� �,��P�b�=�k�}� �ρϓ��Ϸ������� ���^�5�Gߔ�k�}� �ߡ߳��������H� �1�C�U�g�y���A� ������ ��D�/�h� S�����yϧ���� ����R);M _q����� �%7�[m ����/}�&// J/5/G/�/k/�/�/�/���$DCS_C�FG 5��}��!��dMC:\� �L%04d.CS�V�/�#=��A VK3CHS0z��/p#>^?�?�  ����2�1�?�7� �`iMU���(�RC_OUT -6�%�!��/��!_FSI ?~I �9 #8AOSOeO�O�O�O�O �O�O�O�O__+_=_ f_a_s_�_�_�_�_�_ �_�_oo>o9oKo]o �o�o�o�o�o�o�o�o #5^Yk} �������� 6�1�C�U�~�y����� Ə��ӏ��	��-� V�Q�c�u��������� ����.�)�;�M� v�q���������˯ݯ ���%�N�I�[�m� ��������޿ٿ��� &�!�3�E�n�i�{ύ� �ϱ����������� F�A�S�eߎ߉ߛ߭� ����������+�=� f�a�s������� ������>�9�K�]� ���������������� #5^Yk} ������� 61CU~y�� ����/	//-/ V/Q/c/u/�/�/�/�/ �/�/�/?.?)?;?M? v?q?�?�?�?�?�?�? OOO%ONOIO[OmO �O�O�O�O�O�O�O�O &_!_3_E_n_i_{_�_ �_�_�_�_�_�_oo FoAoSoeo�o�o�o�o �o�o�o�o+= fas����� ����>�9�K�]� ��������Ώɏۏ� ��#�5�^�Y�k�}� ������ş����� 6�1�C�U�~�y����� Ư��ӯ��	��-� V�Q�c�u��������� ����.�)�;�M� v�qσϕϾϹ����� ���%�N�I�[�m���ߑߣ��$DCS�_C_FSO ?������ P �� ������"�4�]�X� j�|���������� ���5�0�B�T�}�x� ������������ ,UPbt�� �����-( :Lup���� ��/ //$/M/H/ Z/l/�/�/�/�/�/�/ �/�/%? ?2?D?m?h? z?�?�?�?�?�?�?�? 
OOEO@OROdO�O�O �O�O�O�O�O�O__|*_��C_RPI����@_�_�_�_X_���|_�_o0o+o��SG�N 7��r`���3�@06�-JUL-24 �21:58   ���{`4-DEZ-�15 02:02�`C`Ab Hw�=��b(E�a�a5n�`waWU�w���i�ZX�_��o��VERSIO�N jjV�3.3.2�lEF�LOGIC 18~���  	Gh���Ny��]~0rPR�OG_ENB  �5dEs�`~sUL�SE  cu�u�0r_ACCLIM^�v��s��sWRSTJNT�wfra���0qMO�|�a�q/r�INIT 9=z����Yq�t�OPT_SL ?�	;��
 	�R575@ch�74jm�6n�7n�50���1��#tNy��*wK�TO  W��o�+v]V"�DEX�wdrb�C`)�PATH �AjjA\KJ�LTVL411550R01\ p��\ RG4\k�G�LISH\���H�CP_CLNTI�D ?vEs �Go ǟ��IAG_GRP 2>����R�C` �	 E�  F�,D�E(p �Dx�5j�B�  =��+�B�C�f�T�Ce�EC�� C����G�SCEZX�B�Gm:jf3�62 67890�12345��� � �  A����A�=qA��A�33A��z�A��A���RA���A�ߠ���5j֠Ba�@�  A�`ApX��B�A�C�C�v�`B45l 5e�W�Ba
բ���W{A�ߠ�ߠ�k�����G�Aď�\A��A�Q�7�� �2�7�F�7��U��ߠχ��۠����������?A�ffA�۠�@������ÿտ[�_���Z�U�O�
AUJߠD۠>�8۠2�,O�&�8�J�\ϾV�`��A[��V�k�P۠K
=AE��A?�8��;A2��+�
�Ϸ�P������[������U�x�q�j�}c�\Q�AT۠L��1�C�U�g�y� [���v����Ѧ��-�=�G�I�>8�Q�U�-�8��b�q�7�Ŭ}�-�@wʏ\���p����m@*�Ah�а���<�C�<�t��=�P=�hs�=�ᗍP-�;���
��<#�5l�Ð�?+ƨC��  <(�U�b� 4����A�����M�5iA@Ab? 5����r������ :�������5Y<kM	?Tz�
�d�-��J�G�-� 2��C`�-�xC����}�
���{CEY����ɦZjH��'�p�}��/��Ҧ�ED � E���D�����m�/  8��?��?�:��>���?�ف�����L�-�
zU?�+�-�����z, D lE:p�C`���`�o/���/J�/�"5i�E)���X��O�BIq��/?}/�&??J?5?G?�?D` ����ϧ�?�?�>�?O OD�V��uWO�FO �O�O �rO�O�O�O�O _�O�O_d_v_T_�_ �_6_�_�_�_o�_*o <o�_Ho"o�o�oto�o �oVoHO:% ^I���i����J��>:��6�-� �og�Iw��������� ��	����?�Q��o x��������ҟ���� ���>�)�b�M�_� ���������/�� (�ϯL�7�p�[����� ����ȿ�ٿ���6� !�Zω?�?�?�ϴ��? �����+O=O/�Aߣo e�w��o��]߿��߯� ����+���O�a�?� ���!�k������� �'�����]�o�M�� ��/���g���G��� $J5n�W�� ��	��"Q�C U7�y���Ϗ�� ����-//(f/ Q/�/u/�/�/�/�/�/ �/�/,??P?;?t?_? �?�?�?�?���?O�? O:O%O^OIO�O�O�O qO�O�O�O�O_�O_ H_wωϛϐ_�_���_ �_��/o/ooSo eo��9o�o�o�o�o�o moo�o+=as �o�Y����� �'��K�]�;����� �C/�_ޏɏ��&� �J�y3�X���}��� ������-��1�/ U�g�y������I�ӯ �ǯ	��ŏB���f� Q���u��������Ͽ ��,��<�b�Mφ� qϪ��?�����ϙ�߀�:�%�^�p߂�LU��$DICT_CONFIG ?m���sVzP�egWS����S�TBF_TTS { LT
����VER��xQ�����MAURST�  LT�՜�M_SW_CF��@���ZP��OCoVIEW��A<�����ώ����� ����XR|��#�5�G� Y�k������������ ��x�1CUg y������ �-?Qcu ������/� )/;/M/_/q/�//�/��/�/�/�/?��PM�5�B<�xS��  ����;SCH �2H<�
�yQ�Schedul�e 1 LW ���R䑏9ZP?�?M�HA8�1�?L[=A�4>L�Ͳ2D �?�?�?O"O@OFOXO jO�O�O�O�O�O�O�O �O__0_B_`_f_x_ �_�_�_�_�_�_�_o�TJafeU4ueD5�9m*o �9Dzhg no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x�����@����ҏ�����5=`6�Jeb�t����� ����Ο���	H�V� �)�;�M��?�?���? u�;oMoo����ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ���_o�B�5�G� �7�I�[�m�ߑߣ� ������>����!�3� E�W�i�{������ ��:�����/�A�S� e�w�������S��# 5GYk}��� I����92�?`� r�c��T����ψ ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?��� �?����O(O:OLO ^OpO�O�O�O�O�O�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �&8J\ n�����@ R#�v��?�?�?H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d��?�o ���o�o�o֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tχϘϪϼ� ��������(�:�L� �o���������
�� .�@������ 3. ���6�� ��v�(�:�L�^�p��� ������������  $6HZl~�� ����� 2 D��p�x�ߦ�d߶ ����/"/4/F/ X/k/|/�/�/�/�/�/ �/�/??0?B?T?g? x?�?�?�?�?�?�?�? OO,O��P�O�O�O �O�O�O_ _f��b_ t_�_�����_��_z �V�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��PO8�tO�ODOv� ��������Џ��� �+�<�N�`�r����� ����̟ޟ���'� 8�J�\�n��������� ȯگ쯒O0_b�t��� ������ο�F_�_"�4�F���4��_�_�� �_��:�L�������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ��������^���4� F��V�h�z������� ��������.@ Rdv����� ��*<N` r�����R�� B/T/f/x/�/�/�/�/ �H�??&?�ϒ�c? ��T?�,���?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_>���_/ &/�o(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z���2/�/ ��&�8�J�\�n���@�/(?ԟ�`�5n� @?R?C�v?4��_�_�_ h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτ��_ ����ԏ揤����� ,�>�P�b�t߆ߘ߫� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�򏐟����* <N`��蟢��  �2�V�����ϖ� (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?�� ��x?�������?�?�? �?�?O"O4OFOXOkO |O�O�O�O�O�O�O�O __0_B_T_g_x_�_ �_�_�_�_�_�_oo ,o��p�o�o�o�o�o �o ��bt� �6����� z?�?V?��,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$��?PoX�to�oDo ������̯ޯ��� &�8�K�\�n������� ��ȿڿ����"�4� G�X�j�|ώϠϲ��� ������ߒo0�ߔ� �߸������� �F� B�T�f�������� Z�l�6���������� "�4�F�X�j�|����� ����������0 BTfx���� ��~�0�T�f�$� Vhz����� ��//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?r��BOTO fOxO�O�O�O�O&�h�__&_�z7���� �_��t_,��_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |����>�?� O&O�?6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v�������2O �O"�4�F�X�j�|��� ���O(_����`_r_ Cϖ_4����h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r���Я�� ���į����,�>� P�b�t����������� ����(:L^ p�������  $6HZl� ����//*/</N/�`/ƿϢ/�/�/@Z8 N_ �2�#?V�?���� ��H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ ���_����_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L��p/ԏ��� 
��.�@��/�/���� �� ??�6?ԟ�_�_ v_��,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� �_p�Xϔ���d��Ϩ� ����������&�8� K�\�n߀ߒߤ߶��� �������"�4�G�X� j�|���������� �����P��������� ������ f���BTf�*9�/��ҟ��� �Z�l�6��� 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/?~�0�8?T�f� $�v?�?�?�?�?�?�? �?OO+O<ONO`OrO �O�O�O�O�O�O�O_ _'_8_J_\_n_�_�_ �_�_�_�_�_r�bo to�o�o�o�o�o�o& h"4F���� t:?L??���� ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ^?o��4oFo o6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬ�Ro�o"� 4�F�X�j�|ߎߠ��H����� �10��k\�្� �ϟ��������"� �����j�5�G�Y��� }�������������B 1�Ugy� ���������Ͻ� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�߻�OO 1OCOUOgOyO�O�߻O �O�OYK�_o��R_ ��A_�_e_w_�_�_ �_�_�_*o�_ooro =oOoao�o�o�o�o �o�o�oJ'9� ]��?�?�?�?�?� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E��?�?�Oͯ߯ ���'�9�K��O{������a��$DPM�_SIM 2I����ʱt������C&]Y&Um� � 0�� DϨ�q���RC_CFG Jʵ�!�X� &]���ϸ������ ��5�6ᾰSBL_FAULT K���s�O�GPMSK � &Tb׾�TDI_AG Lʷհ�SQ��UD1�: 678901�2345��xz޻P �����1�C�U�g� y������������X	��Y�۽@��ORECP�ߪ�
�� ~�ܿ�ߴ���������  2DVhz��������9�K�U�MP_OPTIO1N|�[�TR��}�z_�1PMES;�J�UTY_TEM�P  È�33BȱЅ�A�o�UNIT|ׅ��Y�N_BRK Mlʹg�EDðZE|��'t�c�x�TA�T��EMGDI��[��NC#1Nʻ ��X/K/&^u�&[d���/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>COUOgOyO �I�!�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo �J<OFoXojo|o�O�o �o�o�o�o�o0 BTfx���� �����4o>�P� b�t��o������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �,��H�Z�l���|� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
�$�6�@� R�d�ϐ��ϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��.�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������&�0 BTf����� ���,>P bt������ �/(/:/L/^/x j/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?/O 2ODOVOp/�/�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_O O*o<oNo`o zO�o�o�o�o�o�o�o &8J\n� ������foo "�4�F�X�ro|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� j�t���������ί� ���(�:�L�^�p� ��������ʿܿ�� ��$�6�H�b�X�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ������ ���.�@� ��l�v������� ������*�<�N�`� r��������������� 
�&8Jd�n� ������� "4FXj|�� ����//0/ B/\f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �OO(O:OT/FOpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�?�_o o 2oLO^Ohozo�o�o�o �o�o�o�o
.@ Rdv����� �_�_��*�<�Vo`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟB����� "�4�N�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�F�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������ � �$�>�4�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
��H� Rdv����� ��*<N` r��������� //&/@J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?��?�?OO8/ BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�?�_ �_oo0O"oLo^opo �o�o�o�o�o�o�o  $6HZl~� ���_����(o :oD�V�h�z������� ԏ���
��.�@� R�d�v��������� �����2�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� �����Пڿ���� *�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮�ȿ �������"�,�>�P� b�t��������� ����(�:�L�^�p� �������߮�����  �6HZl~� ������  2DVhz����� �$ENETM�ODE 1O��  
����������RROR_PRO/G %�%��:/�G)%TABLE  �%�/�/�/��'"SEV_NU�M �  ���� !_AU�TO_ENB  q%�$_NO�!� P���"�  *�20�20�20�20� +10K?]?o?4HIS�#����;_ALM 1Q.� ���2<��+p?�?�?O"O4O�FOt?_OUT_P�UT 2R�= G @ٌ7���$_�".0  �01���J�TCP_VE/R !�!2/VO�$EXTLOG_7REQ�6�9S�SIZ_TSTK�;Y 5�RTOoL  ��Dz�2��A T_BW�D�@xP�&�Q-W_D�I�Q S�4�����VSTE�P�_�_��POP_�DO]_�FACTORY_TUN�7�d%iDR_GRP� 1T�  �d 	�O|o�m`��[���.���FT&�hB�( ����fmc�o�mm`�C��C?A}�C��B���B�ٙB�$��mArA���AA���Aj��A7e�A�� ~�ٸ�o�oK�qr��HB|���B}A̩�#A�ffA����m��l�E����QW5���\��+�����K�m<��><�`�ws��
 G�r�Dq�q��B����2_q�LZO��:�s��l��N��B��ƈ���m@UU�U��UU\�叀� �E�� F@�����mOHcG�P8�L�u�S@�K�y
�m?x�\���:G:����9{�����m���8����?`�q+ �4��9?����T�ԏ�o�o00%U6�j	��o 0�ۏT�?�x�c����� ��ү�������>� �;�t�#���9����� ڿſ���"���X� C�|�gϠϋ��ϯ��� �����͟?���� ��%߇��߫������ ��,��P�b�M��q� ��Y���}������ :�%�^�I�[������ ������ ��$6! ZE~-ߟQ�c�u� s�o D/h S������� 
/��./@/���v/a/ �/�/�/�/�/�/�/? ?<?'?`?r?]?�?�?�?�?�?\JFEAT?URE U�U�P�	aHan�dlingToo�l 'E�A�E�nglish D�ictionar�y-GMulti �Language (GRMN)0D�4D St@ar�d'F/EAnalo�g I/OzG�Gg�le Shift��Outo Sof�tware Up�date�Imat�ic Backu�p+I�Agroun?d Edit @-G�Camera�@F��OCnrRndI�m�C%\ommon� calib U�I SHVnQSPMo�nitor`[tr~%@Reliab�@�,HData Ac�quisoS�Yia�gnos�A�A*JD�ocument �Viewe{R�Wu�al Check Safety[Q�0Fhanced �Us�PFrP.Gxt. DIO kPsfi�T(gend`ErrzPL�RDmg�sCir�@3` BW�D*JFCTN M�enu`v�S�gT�P In�`fac��eKEG Pp Ma?sk Exc`_@�KEHT�`Prox�y Sv�T�fig�h-Spe`Sk�i;T�e�P7`mmuwnic�@ons"x�ur�`�`=_�A�bc�onnect 2�Yxncr�`str�uAB+IKAREL� Cmd.XG�{R�un-Ti$`Enyv�x�`el +�@�s�@S/W-GLicense�S�\Z`�Book(Sys�tem)*JMAC�ROs,r/Of'fse�@LEH7`�@�J�LEechStoEp�atpp�RLEiUb��Kt�x`�@�@O�o}d�@witch���opR�Q.E�ȋOp�tmڏЃ�`fil��\τ�@gOwLI-T��`
S+IPCM f�un�wP�o�TRe�gi�r=pS�ri��PF`����@Num� Sell���"` Adju-p��ϑ�J��tatu�����Z�KERDM Rob�ot>@scoveLGA4�emj�7anqG|4�@�Servo7`���,HSNPX bx�r�N�CLibrFCD��@ {�����o�p=t�`ssagI�0DTCP �C8�)K���/I�m��MILI�B!���P Fir�m�B�P�cAcc<P	[TPTXJ���eln8�>���$A4���orqu�@imGulayQQ��u���Pa�q� P�Qփ&��`ev.0DUSB� port SPi�PN`a�P,�nexOcept`Y�n�SX,�h'MVCWQr8r/rp�V�P��\��ű����SP CSUI�����XC)KWeb Pl��y�O-Ԁ�`d�Qzf?��f�G�ridD�playP`���Dz�R��.qJ��ۍ�AAVMuyd3epNa�PAxy`Xy�����R-20�00iB/185=L|Mscii�aΒ�Load�P\�Up�lr�Oto���`opPBA�F�qW���(Y�E�`rk��QPR�UT��SRT/K�eybowAMant^@v�C�Pl sd��by E-c�HVl�:@qQGuwF<�N�PT�@cXss@t �t���HV�prE�s@�fUyqc�@�r��ori`>�VCS Jo��s�c`���a�Blu�UH������Pmain )N#ay�.�Yy���N��ifi�SmDG@�p+JUb�Outp�uͲ(g���imiyz��KfAxis7a��Q|mm��s���fR�L �"`��eMI 7Dev�p (���fxvteΐV�PM�X�b��^�/C֐o.F	J��x�o��z;�H�dЃ.FO���Qb��P��oS�ROFIN�ET�J�d�GR�AM/JOG O�J����FPassw�ol�i��񸍇��`C�li�Q�P��EE?D OUTP��d��`�d��s=kVAG�n�rx�� `vog�i 7��B�*��3:�e#avI��ߋ�V�KE?64MB D <?�j3FROs;  퀉@rcҐvis�zS*D trs�Ax�x�.@r
!Pe�ll�L.@INT &MVsh�1(Fa�`�<=c��AD p�7�@}p� " #1�7�ty�@�  x_�lo����(rsv�\��� � p1`�Sd8�p��w�./s��PR(D�� 2P��Q7�� 
PCV`MAsILR�6 e4.,@�E% �Pu+ fx_�mh?�x��Pq \̺2fT1G�Tro�du�w40� �� �LOAD�s  c
P�``�,��4�S[�.�PT��p^u9
! n�SN`N�`cro�`U��� �p�Syn.�(RSS) PR{INU�quiry`		 Zq�����(Ds�\
�QestDDSm0�t-  \et�PS1S�) ՠteHP�nom,@S7@��m�iLj-fle��px�a_�v8H549�$�r'�dib��d��P1 cR��)CTrp�|� FE@�d71{apa�9�Ub	P�#{aZ�Pu}ie�stdpn���S�@�#V8.x pI�\T�!EMZ$��EQ ñ��END�IFREU ��e��d%a1  .�@�s\0� +ޜ0ete"}�wh�en arg��f�i��͡CD�ti~8*.pc pA'�͡u8d R.S�kif�WF,� B�CK 8Ab�v�q�ung�05��!r�
�P�!1�1%��Q�A� F�`b.Tig�/T�ix up��� l�bof G=O4�To f��G��p��mN�F�s��tQ�3�D-PS-�s�rj�Diff.�a.d S.PN:?FW-CHK��
��CD:��SST;EP̢BWDk����.Er.af� 8xVag_C+��sseJ�� Iss�8`�+P.Allo?c.Mem.쀛�k���m I��w .�K[�l Var.�Scr�����FBw_CMB�lar��܉�I�wr.�!FUNC-MP�-���	p��R�˓k�n.sMP�8Z�cmd.e;r.-Pdl.�Pהx��b�'SignǱ��&x�TSHELL� Hepbeat�8No�.On}/��w.SRV��Ў��,�9�m�� a�w��GunM.D�O.@!.Gen.��A��?�.scrn� freezG��P381+Invn9`ig.��ch��x ABC&"gj��'!.d��.uP�p�.��aו4�.��.�abd PGPXtk�k�.��spdd�ѐ4�  k|���0�� pcls<��۳ripcտ��BQ���B�/�no�pa)�K�hgri E�g��aσ�yR~ϟ��mhse�ϻ�\m�hg����)B��̴I
����v	�+�t���%�G�^P A�7�.v�r]��!�1zߛ�l �߷�q����q�������$���^Q�'�"FCT!���_�UrZ�{��CVLOu�k�rcy.���val\����B�����ߪ�r_w��U�9�s�w�2zPCq�7�_tp�N�`�AP��ϝ�wt�� ������W*@x߂��_pr��F���70$�~R��e����sTX��f�"SI1&Ssi��of� i�;�s�G H5<��SPLG�g�gII)�˴lu����al����@-/S��RDEI/k#760H/�$P���/�} �/��������t�@�/`ptk?�ĵ )?K31.�E?��e d/�4��P<�r?�>�	��?��t\j�?��/@�/�&��%O!r�NE576�Dj�0�F�0�/f�He`���0P/p_��th��6�!j���{^��Au_�γ]bwd�O�TER9 �f�RBW�_'�9R o��P9og� �! _f�-�_Y/�o"8�Щog�Lib�ok�}_�_E1?��V
IFpo��D_����#\a8�j_�~1��D�m4RFooE Eq�1��D870��U (̌o�EI)h���d2x4FߎNDIFُ��63.f���o���63��2��k�w2�t/&�Xj8�g 9J��ۓ) "`?��'utx�w$2��͏�J�!O�/��;�2t�v9cO��j72���?p�O_��*�vrc�G�2\w���?�on���ﵿ .�P��ӳ�[Ϳ�`@OB9F��^yrs!����e�/�V�Y���mp��_�5DE ��O�, $�n�<�����.��IߣT]09�/�it̿�41���F�/���06 H����H6s29��w$ H7�߆�12�ߞ�Я;�9�9����63Q�s�M�T (m���Q�FS���mt(�� �U�t�O�F8�ߒ%os ����M��dsg���N�� Ax��T��@�����g�0' x�&��F �kg��e̛��de���! ��o��o��X\O��din#$��l��o��R��WnvL��-���FLX�Kd� �4x_��*/���_`/  870��%)� y/��u �//e[/If5`8�/��=ion�&� 4�F�g����Y?O6��$�4^�r�?�3Fm`�?�$M-1�?�5 d�?G�0_Ŧcl�� ��y�UO/�ɰqO��si_\��Dj59�/ �DB��?/,/>/��9_g 02��=_n�O��\w�?�OLv��o��_\�
ojO;ngx/ƥexXϚ_�_�_  ��P�os��.dO_���d�oƦ50�*UfdL4_R%pl��EJ+��m��/I/��-Gm ��oo.o7t�oK��! i ��%?��oAa|��B���\_�0A�Pя+TvrH�e ]�	�s�������~�͏�_��;�E��4sd@��v>�P�%�Ha,!� �$�@=��)��u���_Z� J���"S�o#���P��[�S" #U�w�Fp �N��h fl_��2q�L���dTo��j�T���%1P  �H552�c�21.� srs�3"���R78"��Q��0W ushJ�614�Q�A�TUP'q88Y�5S45/SY�6[�jp��VCAMo�! �CRI�� - �E��UIFk�ni�fY�28ã��NR�EK� R6A�63x.�~pp�RSCHs �8 JDOC�V����CSU  �R659Y�0^�e�t SEIO1CG�q0A�54"������9���A�SETΣ�csnq���#1�
Y�7���@d�MASK��\h�(�PRXY��DI�F��7��z�OC�OK�3.1�3o0l�ibq�"�MCal�1�R�� ��J6Q�6;69|�539����� (iRL�CHN�1OPLGo3q�0~Т�@��MHCRG�MCSj�mg���Ђ�q�q�y5��%�MDSW�Pmg_�q����q��!�MPRr�g_ex��f�a��R��P��PCM����x���Q����f�ju�1�v�51pf��A��v�3\v�GPRS*��aY�9fоU�FRD��rwecpA�MCN_��H93R�Z���SNsBAǓ��HLB{�{SM��! cv��^��Visiq�2R���p��HTCj��!_TMIL��6���C���90��TPA�� R81A�TX���L��TEL��V�T (�Ү�CP (�J8E���C�.�=ÇJ95��]��f�i;ni�UECN�a�wUFR��\cv��VCC��B�(�VC�O��� ��IP.�!����SUI��P�C�SX�t (��W�EBj�
_�HT�Tj�576|�R6�2����CG (�ABIG��(���IPGS�% R�C.���P�88��t�\r5�89v�i� "P�W��W��H]6}�ui.�7ш�0|�x�
����d������� Px�6�1����< J8��JC89����v�V�aq��7�� (< R53���� ��68��y�66��R74��L��~�ps��5v���q��6��%�R5ti-b4�J7% 9�A�l�ѕ�98v�6\��e�]�82��Eq1Ң�r.��56VMo��65.��55^~�R DM=�6R��H7��5��99 H��6�� ��"�U���.�DRc�6Yo;r d�R64.�9�J��E9��t\d�m���� d�s�.�
�EN(!69~ЉR=6��j932�����sit�98��or������П�j!�INT��~����5>o0���du������� D06��QA���"pstr������SVMrй�CLIr�tr_H��v�=ÇCMS�I�� j�_;dcL STY.��p����Z���CTOj��n�`����Q9�3�2$�JNN��y�N�N��ORS��2\]p4�R68R�c�"8s���"EXT6 �#9F�ҭ�OPI6 ���S2 �"l2!!�$PRmQG�RL��_w��Sd257f�!3ETuS�1y/1SLM*а����Й52����*0)�CP��2΢�TOA��TR�AN�%�FVA��t;mg� IPN.�=øH@.�I�EZE�0i�n/1UPD~�93PkMC~�8F2P1I�fu3E0��400"�vtm�C~�=Û@��
eD0��sNP�B��}D	1��E7bA�Efе#RT2�Bp� �@���)�@��5�P2QqpuL E0�ѩ�7P�.�m���P~��@T�28}��P� P22��)@�)Q��u3sP�H}�vt�vqqR����P24p�!��7P��mof�R�4��]�S3U�}P27v�58��P���T��7Pv�ER��P3����P4�1�U�5�v�dQ5iQ��|Q�5I��P33~�zvsy��9���E���\mnu=e��������sy� ���be �ne��eް=e���"4=e���4��=eްc=e����=����0�felp.=eq����r�hQ2�e^1�e\i�f���5.utfl =e)���5���k��=eM���Q 7=eqB��92@���`�vR0HoZai�`
u��. ���- �Ђ��f��oK�? =e0�>�eJ91=e90i1�f��9�g30=e�13c�R7p�73�8�fz �gU�=ene^wgisn,=e)��E��rc�vAy%��o�Bin]w��e��\���v909�fnE�=eg�!�e����!���bpfk=o[0j9������f��lf VGqF�f&���J90���2��68��6868�f���J84��y"���ivn���u
��e|ю pvgf�f<N�� gfs�����v1"����s�/�V�vCCR\���r��ڵ�56�90�f46��w�Фv(��fRG�J|crg�v��{F'�rg� ����gxf�ٿǵu��yq;�%�  ��zQ�edfG�Re�jur ��O II)!{�4p�\.0ؗ! jA�!ٟw�ck�vF%�]x4�*R�g݇u�fn���fة ���et�fK"c #�o+�ivguH�0I�!�o�� (lff�p,v�ov��erv ���Vej65����aR�6�3\�v�Wdvwe]w��"�5 ����+mz vFr�6���@�f�r,v�P�4�P�vtu�v����AGa ��q��th_�f:�{j��_vwp� �I��� -%�p 2`� y ��c�sexf�9>�P�au ��6E5��u�Ϭ��3� n ��j�����u���T�p��8�6\�v�Wd�sh4�g}ber_���O�w���f�	 �J8̗jo�o2b����R���R����lt��w���� �� fv��f	�h�M� G@A�5<P�oftw�v} 8��0� "F�}���cm,vF`���wal �6�p�1ag��OENU"=/O-MvLi/{dkp�/�.n4朱/�/ARD�/N.P��?�m��)?�%t�xfM?_?PPLt:�  H55�@�#fl!I  �1K !I (M�-!I9!QJ��!Ic3� "!IP=P!I74�\pQJ��!I�Q�K.ްJh774�Jd.�f!ICQ�!I832t�J�� QJiC,!I<!a!I\ngh!I�1!Ig�@!Ir�P!IQ��!I3B !I��H!ZC1,0Z�1�[dr�O�H@�P!I�P0ZM�!I0� .qZ H7!I5��!I:�0O�J10\!I�� 1j�\��!o#GE�Ao3h�L�_�K1pZ�M11<o!I-30i!IM8aZ��Az500QJq�x!IA!Ib\p5�[EN�k�[Z�PZI��[�PRQJH68QjP��o!Ip70�O2ip�/�_X4�_!I/1�5@_RY=�a_�H0a��Zs�\5S���6�J��!ZA/{�!It���0�J! pPj=�m!I>��zN �Z�Ѐ�Zm�Pz~ 0Z51A�PPji�k @�ΐ�J%�v!� "�Z(P-Pj ��Qz�a�0Z��oXq-/K]o|fleъ��0�Jt\`ZAC"80Z%�J "C�3h�\c�|TXaJ\hd��#�C�C31�̂�QZc40JM^h8a2я#G��CS�ZtA�q�j �r R��[ J�m���|@� �Ѐ���Q��Yp��e��ʡ��c�� �O��hs�Kj72 �83�Kn BPz=�Ѻܥ�!IJ78��Biqn0ZmOKact�<� @�ikavA��X�\ikZV�J83�jaQZj7���p��"�4��m�K��npsos��#Gkin�Z��liGE�"�-� "�=�"�M�"�]�"�m� "�}��~�"���"��B�"�oN�"����ko8@���"�prw 
�"�ik�"�4�F�X��j�|�������2ni����
ial��2s'chn#	s = Oas�
�4y���`����B�oc��4�n�3�94�@�D OU�=��M�.�(TC�T^a�<mb�694\�mRx����p "T��r�4\t�*-��z=�5�Spee�L}��24�P�) ���NM��*M �icti�*N���)N,v�/rr�Int :���*��N�RS1�*ce V�*��:��K��r8.pd!Iw�J��rmm!*<��r8\hi0!I>�A!I39\n!IE��?M-�*�0p*��0�*27 (�:a9r��Ngnk�:�� �J�Z��).��N\r�0h�:n\/0.�*@���)��RI=��:)?;��-"M0�*�)f�m�J��r8}�BOt68^L>p-�K���9��r8�H81 *-_�Lm14�*]_8�*13[�P�*741.�*}�A|�.��*3S�2).��r8hMp�:N��d8G �:�NM`QJ.O�Z-O��
E�:fdo; G- M�?�?Ew2����o�l2s�I74f!�CM_:sl�* =⒋�*-�?����+^|�-2/��9͠a;Lo!�M��oo%g_�2o�DipZM�_�q���Ew4�����ĉ�Zݏ�44�/}�70O{A(B�pZ����3`:}��m3�𚭯7�J���[36a ��@�¿d�v����3���o�l70 *2�03)�KTX!� g�Q�s(29P�^/p+29�pp?�)SH6pZ�?h�0�\-/?,M-9!�>������m92��~63�JP� !���9� �υ�90�J�O[9�3[��a�ʮL93q\ ��*�H79 *z�_7`�iB/7*`�P�*�P�II`�N�]7 "@��-5�p���C��o�jL^}96p��B/4 �n?�G9B4@;��b��`�O�N`�M���37��DM�L7o��C�3�� ���-�?�Q�pZ=�?]czla���`�98Ϯn`�799�/1pZ����2�n��j��@Jdz�m-��/�d�n�1750:�P��P`:000`;� ���=�9N���m-�m0H.��H61�Jd}p�1B oҟD'R20oBjAr�"�4��-1���~pH  �STD��15LANG�#1E�q%E�h611%E21U�"%E=�%E\Q@%E ���%E  �%Ew�[yF- V%EOaini%E}�I%E�CVSU%E12 �JyFR68%E68�6HF�@9%EJ84q0%E-�%Eg C�F�on VUIF,�%E~0yF�P%Eetu\%EVI�G]�%E�t\cv%Elmn�HF�%E��%Eu\v!p%E-��_�Rl%E �FuVu.f%Ej5�12%Ene+W. 
vyFJ5TF945HF�0�X� naFine�V��%E��V�Ylnql@fM!yF! j�H1!%E}�!Vst�F�uR�G8TF021DV���dyF(i�fic�s8_J\iag\VIRDG%E��V0�Fw09.�Ve Cf:x09 �h�G�mx�(QVck J\9\�ssiVC"HFEIj`Qp%E�1I�et�v� SS�Vtext��v��F51�W R�7	V683R�BT��I tP_�N�]�ETSS]�r�rorOPTANkӍ�������e��sspc�������Ȏ��bʅ-W`��ce1�����90wpʅJ94�&a��M���
�9)�3�@��q����641��erfa�Ɇ:B��EB��pciMf��v.���pՏ�  0��lވ�I`���P�]1��td��dy���i����r.��ȭ1��@l/���st8S����0 H0@��!�enk2DPN)@IFǁ����N��527����8��෣����!���ene ��ơ!�	�b
��b� ���6�
�A�����b¥(AD�rVa
���ܐ�ARC��7�4���!	�v\aw	�VS�p
�������d��±DǺP�awg��
! o	�~�ئn�s�����1�0@CU�Sa��ܐgí�e�T T�g��e�qRf���b�e� RRESe�5B�f�1�6e�3J9�pf�30K���\�g�692|�22�<g�y�b Pl��:B8Ӆ��web���#htW�ӺPCՍ1��s\hx��R�l7us.��vcp���ame��cՏ�CA�M|ƍ��H558R��L_p��8�9�@������@d�up��R7]3��3 ��C��nE�J88P�47`x���!E�(CamE�B~ rE�mE�0tE�mnP��ł������O\etcE�ư#���� ��a��>���alCib��:q��N H��GH57E���D�L�����2�45�2g�y�o��b UI�}0E�<]���uif\E�5P�E�9r��1E�iew�.E�gr��� J�695��E�6J�4�P�74'�q�R�694�m Vt���qR��t\t��pvw4D� Empvt�ΐ8D�����Dia����MDCR76rL�4᠁�R71E� �`�q��@� E�~���b`Xe�v�:d\���GPT<����nyd�P�skmgE�7cke��ngc��� �b��A�%3'��6�49��ON��c��$83wp
��6�i8N�0�1 4&�`3E�>��J� ���"Ѧ@,�a`��.s@tphE�M������ �.Α�4��J�)� �@r%� �81XP�B�(�S0&5a��A��a��(T��agq.����dtr��,����sf|�R�(�m�	G 	G uE��T�EME�����$	F�E�����&ST�E�?�M�p&>�(���5% q&�Q
Ex�O+ 16��HCHt4&ijHp "�62j�V�?[�s.�����I�pT616�tcpTCP/`��� �^�1�	�~@@) l!  LNk9NB�$��E�W�� OE� ��X6&1?�& L'62f55�Z&%�^��54X&0i`)/�B&�6#8FkP�90�g6J)6;7���h����נB&SX&��2l�/8R7P�68'o9 PTQ�98 e�w�TC�6n�h��v�$pi��"HC\v���%u �wp�	\v��,F�)G�(��k�^/ hcp�Eұ�FX&ry��ʡn6eh:�NmionV�f_�,E�)� �6��:��p�wCTC<j T6\aP�H0�?�4U�@�6�0ݏ��&PL����p�6g'W�)z��Pcri|����tc{��ost���E�F O�g! �C獢"wP��2 )�T�TTP��@�E�_T nE� $8F$V�WEC �/^!�iPR\55����R�NNf38�jp&7B蕪RS,wj9��Ew
?�6��JA�iv��
O_ �^�e�!�@�f�����AF���=�E�}������0����|�H:P�R f0\PR�99��>_���$FEAT_DE�MO U����3�;�p�  ޸N�D�Vσ�zόϹ� ������������I� @�R��v߈ߵ߬߾� ��������E�<�N� {�r��������� ��
��A�8�J�w�n� �������������� =4Fsj|� �����9 0Bofx��� ����/5/,/>/ k/b/t/�/�/�/�/�/ �/�/?1?(?:?g?^? p?�?�?�?�?�?�?�?  O-O$O6OcOZOlO�O �O�O�O�O�O�O�O)_  _2___V_h_�_�_�_ �_�_�_�_�_%oo.o [oRodo�o�o�o�o�o �o�o�o!*WN `������� ���&�S�J�\��� ��������ȏ��� �"�O�F�X���|��� ����ğޟ���� K�B�T���x������� ��گ����G�>� P�}�t���������ֿ ����C�:�L�y� pςϯϦϸ�����	�  ��?�6�H�u�l�~� �ߢߴ��������� ;�2�D�q�h�z��� ���������
�7�.� @�m�d�v��������� ������3*<i `r������ �/&8e\n �������� +/"/4/a/X/j/�/�/ �/�/�/�/�/�/'?? 0?]?T?f?�?�?�?�? �?�?�?�?#OO,OYO PObO�O�O�O�O�O�O �O�O__(_U_L_^_ �_�_�_�_�_�_�_�_ oo$oQoHoZo�o~o �o�o�o�o�o�o  MDV�z�� �����
��I� @�R��v�������ُ Џ����E�<�N� {�r�������՟̟ޟ ���A�8�J�w�n� ������ѯȯگ��� �=�4�F�s�j�|��� ��ͿĿֿ����9� 0�B�o�f�xϒϜ��� ���������5�,�>� k�b�tߎߘ��߼��� �����1�(�:�g�^� p������������  �-�$�6�c�Z�l��� ��������������)  2_Vh��� �����%. [Rd~���� ���!//*/W/N/ `/z/�/�/�/�/�/�/ �/??&?S?J?\?v? �?�?�?�?�?�?�?O O"OOOFOXOrO|O�O �O�O�O�O�O___ K_B_T_n_x_�_�_�_ �_�_�_oooGo>o Pojoto�o�o�o�o�o �oC:Lf p������	�  ��?�6�H�b�l��� ����ϏƏ؏���� ;�2�D�^�h������� ˟ԟ���
�7�.� @�Z�d�������ǯ�� Я�����3�*�<�V� `�������ÿ��̿�� ��/�&�8�R�\ω� �ϒϿ϶��������� +�"�4�N�X߅�|ߎ� �߲���������'�� 0�J�T��x���� ��������#��,�F� P�}�t����������� ����(BLy p������� $>Hul~ ������//  /:/D/q/h/z/�/�/ �/�/�/�/?
??6? @?m?d?v?�?�?�?�?��?�?OO2M  )HHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0�  1�,�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿@޿���&�7�:�-�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�?��?�?�?OO&O8I��$FEAT_DEMOIN  =D��h@�3@PDI�NDEX]KlA��P@ILECOMP V����A�kBKE�@SETUP2 W�E��B�  N� �A�C_AP2B�CK 1X�I � �)MAK�RO900.TP:G_3@%�E_?Z!&_c_:G�E1__�UT1]_C_�_�_y\2�_�_UT2�_�_1ono"y\3ooUT3eoKo �o�oyU9H�lJ3@�@8u�( ��^���)�� M��q������6�ˏ Z�ď���%���6�[� �������D�ٟh� �����3�W��P� �����@�¯�v�� ��/�A�Яe������� *���N��r�ܿϨ� =�̿N�s�ϗ�&ϻ� ��\��π��'߶�K� ��o���hߥ�4���X� ���ߎ�#��G�Y��� }����B���f�����1��K�@P�O� 2�@*.VR:���RP*����#S0����yUn�PC���RQFR6:��4��X��T|@|��y�_@I�xV*#.Fq�%Q	��<�`�STM� ���" ���RPiPenda�nt Panel��H�/�/�8Pi/�
GIFs/�/���/F/X/�/�
JPG�/!?�?�/�/q?F��JS{?�?RP73��?O?%
Java?Script�?�/�CS�?(O�O�? �%Cascad�ing Styl�e Sheets�TO~P
ARGNA�ME.DT�O�l�\�OUO�1�D�O�O	PANEL1�O2_%�_[_��_2P_�_EW�_a_s_oZ3�_:oEW(o�_�_�oZ4Xo�oEW�o�io{o�DSHEsLLp�A %+r�Cm���GZG?_MENUE0-O��u�q���EEI�NGAB�J�%�3�K�L�����vSU�MM_VAG.D$>?�O:���������yTPE_STAT:��;�S�y������E;�INS.XM�[ҏ�@���o�aCu�stom Too�lbar ��yPA?SSWORD�oU�?FRS:\C��� %Passw�ord Conf�ig���G�CONF1��]��Aǯ�����,��yEXTSERVOC�U�K�c��������UIO_SET|��%�AϿ	����4ϣyVWEMZROUS�e�S�kϑ�ؗϼ�K�AGV�UP [�m����ϙ��@��� d�߈ߚ����M��� �߃���<�N���r� ��%����[���� �&���J���n���� ��3�����i�����" ��/X��|�� A�e��0� Tf���=� �s/�,/>/�b/ ��/�/'/�/K/�/�/ �/?�/:?�/G?p?�/ �?#?�?�?Y?�?}?O $O�?HO�?lO~OO�O 1O�OUO�O�O�O _�O D_V_�Oz_	_�_�_?_ �_c_�_
o�_.o�_Ro �__o�oo�o;o�o�o qo�o*<�o`�o ��%�I�m� ��8��\�n���� !���ȏW��{��"���$FILE_D~�� 1X������ �( �)
SUMMARY.DG#�N�MD:W���s��Diag Su�mmary����
��SLOG��p����۟�����sol�e lo����TPOACCN�v�%^������TP Accountin=����FR6:IPKDMP.ZI
��j�
� �����Exception$��ի��MEMCHECCK��������/��Memory D�ata���� ��)��HADO�W������)ϸ�S�hadow Ch�anges,�ߴ�5)	FTP�Ѓ�χϲ�1�mment TBD���ܷ\+�)ET?HERNET��͎�f���3ߪ�Eth�ernet 3�figuraC�����?DCSVRF�ϊϸ�ϵ߸�%z� �verify asll��cĐL8u�DIFF�ߓߥ�:�%��dif�f<���f�z�CHG�D11��*�� �Q����� |}�2p����C� ��j���GD39� �2���� Y���}��UPDATES.� ��ЋFRS:�\L7�Upd�ates Lis�tL͛PSRBW�LD.CM{ό�7�N0�PS_R?OBOWEL��g�:SMp�)��M���/Emailr��aïcĮ�,�� �Տ���� /��$/ �H/Z/�~//�/�/ C/�/g/�/?�/2?�/ V?�/c?�??�???�? �?u?
O�?.O@O�?dO �?�O�O)O�OMO�OqO �O_�O<_�O`_r__ �_%_�_�_[_�__o &o�_Jo�_no�_{o�o 3o�oWo�o�o�o"�o FX�o|��A �e���0��T� �x������=�ҏ� s����,�>�͏b�� �������K���o�� ���:�ɟ^�p����� #���ʯY��}���� �H�ׯl�������1� ƿU������ ϯ�D� V��z�	Ϟ�-ϫ��� c��χ��.߽�R��πv߈�߬�;�������$FILE_7 P�RF ����������M�DONLY 1X��� 
 � q�H��l��y��k� ��U������ ���D� V���z�	�����?��� c�����.��R�� v��;��q �*<�`�� ��I�m// �8/�\/n/��/!/ �/�/W/�/{/?�/?�F?��VISBCK�#��2�*.VD�M?�?0FR:\�f0ION\DAT�A\�?)20V�ision VD file�?�/O O3?AO+?eO�?vO�O *O�ONO�O�O�O_�O =_�O�Os__�_�_d_ �_\_�_�_o'o�_Ko �_oo�oo�o4o�oXo jo�o�o#5�oY�o }��B�f� ��1��U��������MR2_GRP� 1Y��C�4  B�r�	 �.�ҏ�πE�� F@��������πOHcGP�&�L�uS.�K�y
�?�J����π:G:�r�9{�~��A�  욟��BH̃C��=NƕB�ƈҕ���΄���π@UUU�UU��S�΁�=���=�L��<���=�(H�>C�s>�I�b����:���;%�9޹p�9��:��� 2���V����ܯ� � 9�m�Əd��D����� �����οϊ���:� ��_���nπϹϤ� �������%��5�[� F��jߣߎ���J�\� �߀�!��E�0�U�{� f��"���F������� ��A�,�e�P�u��� ������������+ (a�߂�d� ����'���� ������� ���#//G/2/k/ V/h/�/�/�/�/�/��_CFG Z��T �/5?G?Y?���NO ����F1732�68h?RM_CHKTYP  0��r���00��1O=M�0_MIN�0r�W���0��X���SSB3[��_ �
D�e; C)O8K��TP�_DEF_OW � p���PGIR�COM�0aO��UN�C_SETUP  ��%O�O�O�O���GENOVRD_DO�6}�mEU�THR�6 dUd�T_ENB�O ^PRAVC��\�7�0 ���_�/��_�_|O�_� �_(o�_Lo^o�_mo oo�oyo�o�o�o�o $�oHZ�o~�h�3ydQO�@1b���r��eB�8��^���
��';�.�N���F��F�3G�R�'	���D;s3���Czffr�t >p0��x��g���B���r�	�y���!�&���"�D�F�x��������n�ɏ珑����1\�>�� :�\�^�����˯Ɵ� ���ܯ ��At�V� '�R�t�v���ѿ�ޯ�����OGRSMTkScrY�p�0w�m��x��$HOSTC�21d�y�0��Qa}U@n���1��m17�2.26.29.7230��e��*�<�N�`�n�e�ϒߤ��������� e	c�fg_fanuc ���.�@�R�b��E u���eB���إ���� ����(�s�L�^�p��������9�	ano?nymous���� ��e�w���t ��������=� (:L^����� �����9K] 6/qZ/�~/�/�/�/ q/�/�/? ?C/D? �h?z?�?�?�?�/ /1/3?Og/@OROdO vO�O�/�O�O�O�O�O OQ?_<_N_`_r_�? �?�?�?�__)Ooo &o8oJo�Ono�o�o�o �o�__%_�o"4 F�_�_�_��o��_ �����o�B�T� f�x�����o��ҏ� ���Sew���t� �������Ο��+�� �(�:�L�o���f���য��ʯ?Ώ�ENT� 1e���  sP!a��  �	�F�5�j�-���Q� ��u�������Ͽ0� �T��x�;Ϝ�_�q� �ϕ��Ϲ����>�� �t�7ߘ�[߼���� ������:���^�!� ��E��i����� � ��$���H��l�/�A����e���������Q�UICC0����!�172.26.�29.861 G#���	2�s���!ROUT3ER��!7`~��PCJOG7�!192.�168.0.10�CAMPRT�c5 x1����RT ��%/�N�AME !��!�KJLTVL4�11550R01?RS--KU1��S_CFG 1d��� ��Auto-sta�rted2�FTP=��!T�V��/�� ??1?C?U?��y?�? �?�?�/�?f?�?	OO -O?O��/�/�/�O�? �/�O�O�O __�?6_ H_Z_l_~_�O#_�_�_��_�_�_o�o 	SM<����O�_to �O�o�o�o�o�o�_ (:Loo�o��0������ �2� D��ZC��og�y��� ����Z�ӏ���	�,� -���Q�c�u�����TH C����'�I��4� F�X�j�5�������į ֯��{���0�B�T� f���ß՟��ҿ� ����,�>�	�b�t� �Ϙϻ���O������ �(�s��������ϔ� ߿�������� ���$� 6�H�Z�l����� ������5ߛ�Y�k�D� ��[����������� ����
.Q���d�v����4(_ERR fF*���PDUSIZ  �\ ^w���>~WRD ?�%�:��  �backup�?guest�T�fx��3&SCD�MNGRP 2g�%� ��:�\ kDAK� 	�P01.03 �8�   6�  � �w�A�w�.� �������W; �x���G `�����+-  ʯ  
b #��!.,�6�����; �C#������S/N  + � / n �u{/�����_����M? �? �� �/�7U�S`�S`��d/�!/3/E/2���1?234567&�? ��?�?�?O�?*OO NO9O^O�OoO�O#;�O �O�O�Oy?�?�?F_�O V_|_g_�_�_�_�_�_ �_o�_	oBo�Ofo%o �o__)_;_�o{o �o,)bM�q ���Io���(���_GROU�h*�	-0�	�!�1�cz���B�QU�PD  6���C���TYP��� TTP_AUT�H 1i� <�!iPenda�n������!KAREL:*$�-�?�KCT�d�v��L�VISION SETM�ԟ��\J��ٟ�I�'�� ?�9���]�o���������CTRL j����
 k��FFF9E3�ȯ8�FRS:D�EFAULT2��FANUC W�eb Server2�
�,>۬�����Ŀֿ����WR�_CONFIG ;k� f2���IBGN_CFG� l��2\ �@\ <#�
~�BeH|�C��?4:�~�L�DEV�`���V�� IO m�a�I�EXDAT �n����EXFL�G���T�FIL �o����O�TP pYݮa?���������	MER�CATOR!RE�CO�� "R_AC{HS��ISTW*��V�,�V� "SE�NSP��TX�Q�999�Keine 0�k� h�\%IB�SC����M�4�8�2@�EW�𛩀�TĿLMTN  ���� �b����������J�SBAD��� 7�^�x�T�DL_CPU_+PCQ�\B� ��� AY��[�MI�Nd� =�rT�GN��O�H����рINPT_SI/M_DO������TPMODNTO�L�� ��_PRT�Y����Q�OLNK 1q�@9K�]o���MA�STE����SL?AVE r�b��OZ���UOހ<�CYCLu�$��K�_ASG 1sY� ����aП՗�~���`�$0c�������a�� ����%/0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b?pt?�?�XNUM��z��IPCH?���O_RTRY_CCNQ�I�D�N؁��8�� �Zt��FO�T�S;DT��OLC������$J23_DSP_ENB�0��ь@OBPROqC�C���	JOGI��1ukL�ad8��?�����O�??"��ۯ4_�pQJ_o_ �_�_R_�_�_�_�_��zO�y8!�O-oo )_;_�_�o�o�o�o�o��o&oJ�B1 +oeNaoso�o�� ���(�:�L�^�9���BAc������ ���*�<���`�r� ����q����C����?��BPOSF�OF�K_ANJI_� K��&�RE_�.Av/���/�����KCL_�L��2�?�EYL_OGGIN7��������$LA�NGUAGE �����ENGL�ISH ١�LG�-Bw �S���S�xJ ����B����S��'� ���Z��MC:\RSCH\00\Xﶠ��?ISP x���0��⍊�ߡOC����Dz���AݣOGBOOK yY�����!����X x�	��!�]�x���``͛���ه	ε���>��ϼ̲_B�UFF 1z(A�ϟ��ߞ /� �K�]ߊ߁ߓ��߷� ��������,�#�5�G��Y��}�����DC�S |ؽ =��͑�L���$�6��H�Z���IO 1}"cJO��(����� ����������#3 EWk{���� ���/Cn��ER_ITMhNd ��������/ /,/>/P/b/t/�/�/ �/�/�/�/�/?��q�SEV@�mTYPhN�l?~?�?=��RS�0����B�FL 1~|�@��OO(O:OLO^OLpO�?TP��y[2}��NGNAM]���6ˢ��UPSc�G�I�0c����A_�LOADPROG� %�%UP�024}O��MAXUALRM�ܑ���筥
DR�A_P�R�Dܐ³ڑDPCf�ع�ͪ_$�;Y��P_GRP 2���[ �S�2S�	[1�0�ڐ�o �V#oo oYoK�Go�o so�o�o�o�o�o�o *<`K�gy �������8� #�\�?�Q���}����� ڏ�Ϗ���4��)� j�U���y���ğ��� ӟ���B�-�f�Q� ����������ǯٯ ��>�)�b�t�W��� ���������ݿ�π:�L�/�p�[ϔ�=WD�_LDXDISA��@+;l�MEMO_{AP�@E ?�K
 T����߀�&�8�J�\�n�DPI_SC 1��M��� ���T�Q���߅���� 2��V�h���w�K�� ��������
������ R�d�O���o���-����������*��C_MSTR �,=~ISCD 1��������� �:%^I� m����� /� $//H/3/l/W/i/�/ �/�/�/�/�/?�/? D?/?h?S?�?w?�?�? �?�?�?
O�?.OORO =OvOaO�O�O�O�O�O �O�O__<_'_9_r_ ]_�_�_�_�_�_�_�_ o�_8o#o\oGo�oko��o:MKCFG ��X�ogLT�ARM_�b�X;�b �c��� (t�b_GRP_�DO �X�a����l�<uq�hk������o$MMETP�U��Xs��`	NDSP_CMNT�8�`�Q  �I���q�al�v��POS�CF"��f��RP�M!���STOL {1�X 4@�`<#�
���a�� � ����"�d�F�X� ��|���П��ğ�蟀��<��0�r�\��S�ING_CHK � %�$MODAEQ�c��o�g�i���DEV 	X
	�MC:C��HS�IZE�͚`Ȭ�T�ASK %X
%�$1234567�89 M�_���TR_IG 1���lX%�ܪ��c��Կ���� ˿Ͽ�<����7τ� +Ϩϋ�aϣ��ϗ������/�YP���`���EM_INF� 1�w �`)AT&�FV0E0%ߜ�)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ������H�����D���AL�t�/������ ����߸�����M�  �q������Z����� ����%����[�  �2����h��� ���3�W>{� @�dv��/� //f@/e/�/D/�/ �/�/�/��?�� �a?s?&/�?�/�?v? �/�?�?O�?9OKO�/ oO"?4?F?X?�O|?�O �O6O#_�?G__X_}_�d_�_�nONITO�R=�G ?��  � 	EXEC�1�c�R2�X3�X4��X5�Xp��V7�X8
�X9�c�RkBOd�R Od�ROdbOdbOdb Od%bOd1bOd=bOdIb�Oc2Vh2bh2nh2�zh2�h2�h2�h2��h2�h2�h3Vh3�bh3�R��R_GRP_SV 1�q�� (d�>�fj��_f�?�
���a��I�?_g+�Ze��_�������Y7�_D�@R���PL_NA_ME !>�Y���!Defau�lt Perso�nality (�from FD)� �TRR2hq 1������Y�  	 d���ŏ׏���� �1�C�U�g�y����� ����ӟ���	��˨2��K�]�o������� ��ɯۯ��<:�� )�;�M�_�q������� ��˿ݿ����
�;��P*�g�y� �ϝϯ���������	� �-�?�Q�c�u�D�V� �߽���������)� ;�M�_�q����� �ߚ�����%�7�I� [�m����������������� E�@ E�` E�F�}�<N�d�tl~c��! 8��  ~q� 'EKi� ������//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?-�F? X?j?|?�?�?�?�?�? �?�?�O0OBOTOfO xO�O�O�O�O�O�O�M �_$�=_��a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�oP_ �o�o�o�o�o�o# 5GYk}��� ��o����1�C� U�g�y���������ӏ ���	��-�8N�\ ���j���� ��� ��r �B�8�f�\� n����˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� >?W�i�{ύϟϱ��� ������O�/�A�S� e�w߉ߛ߭߿����� �� _�$_=�O��s� ������������ �'�9�K�]�o����� b����������# 5GYk}��� �����1C Ugy����� ��	//֟8�N/\� ���/���/�/ȟڟ7/ ?��??&?8?V?\? z?���/�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ >�W_i_{_�_�_�_�_ �_�_�_�R_/oAoSo eowo�o�o�o�o�o�o �o ��+6�O�s �������� �'�9�K�]�o����� b��ɏۏ����#� 5�G�Y�k�}������� şן������1�C� U�g�y���������ӯ ���	���/8/J/`� n/���/|����/2��/ ψ?�?�?2�8�J�x��nϜϨ��$MRR�_GRP 1���������  �`� �� ����� �@D�  ��?������?������@T�;g�Ũ���*�;��	l�	 �����X��'���F�O��^ �,X ��k���K��K��CK�zK�~o�K{GK�M�sA�S�������?�;g?���N?Ę	@�
���Р߯��I�ۿ�
���������X���4  ��p7���ô�7���A��  ���Pտ�n���'���������Ѡ���(Ѵ�����������  ���������	'�� � )�I�� �  ����O�:�ÈM�ß�=���e���@u�{�v�����������������������@�?�ɿ@{S�@�@��)��C6�B� ' CaK B�B��Q������C9���L ���� ��}� H��B��� ��0 ����Dz�� O��$J!�3�jnz  ȅ:=y��� ?�ff�ؿ��O ���,68��/(*	�H��=$0(��V%P_(�z��U�UԿ�?33�3��6;��;�QaT;\��;���;�	�<�$D���/�A04�+���?f�� ��!?��?&0��A��5@�, %5�q1�-��]? ��|?�'A���?�?�? �?�?�?OOAOSO>OwO�F5F� fO�O bO�ON?�Or9�O+_�H�E�  E;�E@ E����Oq_ \_�_�_�_�_�_�_�_ o�_7o"o��jo���o�Jo�O�o�����*�G\h�H�����?0���` ?E�jfB�'o �$6�*���?�	��_s���@�������yA� A��t��Uq���7���w�(��|?��`d�k�������ӌ���k��C����`L���h~��~�}�!�� �%�D/�C�G33Ck�B��1B-v�=����%�E��ីW
��u���²B�����pX��Blz��X��}�����
=Õ���ö�=BU(�������F<rѾ��JD��LUW��H�� I%K�Ab!&�LU�L =�L]���HP� H�R�����TF�L%��J�
`H��H���A�� |�j�U���y�����֯ �������0��T�?� x�c�������ҿ���� ���>�)�b�M�_� �σϼϧ�������� �:�%�^�I߂�mߦ� ���ߵ��� ���$�� H�3�l�W�|����� ���������2��/�ph�S���w�G�>���� C��\s��x��Ć�����CV���L7��\]G����(���`����!�y���$rc�<�A3-NQ!3�A��vM_�?�v3�g�y��!�;�%D93ҵ�����	/P�-/,V�P�"P_.Z�{o�/��/�/�/�/�+)�/�/(??�8<�8?G?Z�8"�t a?#?�?�?�?�?�?�/`mo'OOKO9K9QO0[O�OO�KO��O�O�  �e 3� �O�O__9_'_]_kZ  2 E׃�jE�`�W�gBg���r�C��	�pj@��_jϜ��^Gr0 F�� G�� D	�C C�X�_:oY��_@�_zo�o�o�oj?� T�ae�4jjr�1Q�\�
 �o ,>Pbt�� �������:T�{��IuD�YX�Ӏ�2A� @�D�PU�?ϐ]� �� `?�aϔA��XU�Ij��;�	la�\!}�����e�<�0F�����������'��0}� G���?}�h�����ş ���P�����V_�z&'��9�G���k����+UUp�s�=��ͭ���Y�Ϡ(bۯ�Z�&f���G�TY3�>�u0  '  [� e�Z������� )b���ҿ��B�P�� [a-�abCp!��T�@��x�cϜχυ�j\����  �j:v�a�`x#a���
���� R�dۖ��0yߋ�>Ρ'`i���0����쿢>Lס ���A����4��e)a�G�a�*�?fff?[`?&g��σ�"i b�)mv�]���[���L� ��x����5� �Y�D��}�h����������_ F�P����7�� X��*�&��� ����-Q< u`������ N/r;/�_/q/�/ �/4�/�/V/�/�/?(�/7?"?�R�_4�P �Qp?/?�?:(�0�~? �?�?O�? O9O$O]O HO�OlO�O�O�O�O�O �O�O#__G_2_k_V_ h_�_�_�_�_�_�_o �_1oCo.ogoRo�ovo �o�o�o�o�o	�o- Q<u`��� ������;�&� 8�q�\���������ݏ ȏ����7�"�[�F� �j�������ٟğ�� �!��E�0�i�{�f� ����ï���ү��� �A�,�e�P���t��� ��ѿ�ο��+�R7=(�����M�_� I��mϣϑ��ϵ��� ����!��E�3�i�W�(��{ܶ5P%�P����4���B����	� B�-�f�Q��u��� ���������,��P� �߹����������� ������B0R�xf����  2K��*<N `r����� ���/"/A�F/T*
 T/P7�ߓ/�/ �/�/�/�/�/?#?5?�G?Y?k?��t/��{�J��4�� ��~�1 @D�  �1�?��3 � `?x7 �27 A�X�5|���? ;�	l�2��}�KC�0"K> F����?/.�?:&�uO�L> �8�O bO@/�O�O_�O%_] �0@J_XW�x_��A�Й_�X_�_U+�UU�_�_=��� okiS/`�09oGh�R&f]oom�2�	�o6^?u0  '�o�h �_�o_x,�2ZO2��hB Px~ 1@�`�u�aEC���o���o�����R��p&�4�  ��r:$h&Nq~U�2�|j�|�� �в�ċ"�q8�pڏ�>.a�0��1�z2�$�L�">L7a��pA�=���;�����s�2�3�2�p?offf?�p?&ǐ ���t�2�4�y�5 ��8=���D؟q�\� ��������ݯȯ��0��7���Ffp&� s�"������2���� �����3��W�B�T� ��xϱϜ��������� ~_,���S߮�t�ҿ�� ߿������ߔ�
��O�:�s�^���-AfpA������ �����ꈕ�o��?�*� c�N�`����������� ����);&_J �n����� �%I4mX� ������/� 3//0/i/T/�/x/�/ �/�/�/�/?�//?? S?>?w?b?�?�?�?�? �?�?�?OO=O(OaO sO^O�O�O�O�O�O�O _�O _9_$_]_H_�_ l_�_�_�_�_�_�_�_ #ooGo2okoVoho�o �o�o�o�o�o�o1@C.gR�vw(������{�� ���'��7�9�K� ��o�����ɏ���یJ�P��P�Y�� ~O��xT�~�i����� Ɵ���՟����D� /�h�S���w���W�� �=��� �6�$�Z� H�~�l�������ؿƿp��� �.�  2�� T�f�xϊϜϮ����������C�(�:�L��^�p߂ߡ��ߴ�
 �ߔ�������)� ;�M�_�q�������������{J������� �@D�  �?�>� � `?��!���A�X��I�� ;�	l!��}��k�e�%�����F����K�������������=����� =(aL�p�y������������z+v+UU<03=���m�����&f�������u0  '/'(K/�vo/��.���/Z(By �/�. @[ �%[!EC0�_/?[/ 8?#?\?G?EO0�?.�7  �O2:�֮!	
�!�W<�?�?n?� �O$KV18O0:OHJ>��)�M:0�?�O�/��>L��V0A��O�?�O�?O3�!��!�� ?fff?� ?&'PR?C_ O4.�"Q.�M9�}_� �_Va�8_�_�_�_�_ oo=o(oaoso^o�oR]`F� �o�o�o �on_�Y�oK�oo Z�~����� ��5� �Y�D���� R���ԏ2��n�� 1�C�U��Oj�|����`��ӟ�����A� A���'�0��T� ?��E�>�����ï�� �������A�,�e� P������������ο ��+��(�a�Lυ� pϩϔ��ϸ������ '��K�6�o�Zߓ�~� ���ߴ��������5�  �Y�k�V��z��� ����������1��U� @�y�d����������� ����?*cN `������ �);&_J�n �����/�%/ /I/4/m/X/�/�/�/��/�/�/�'(y����?;	???-?c? Q?�?u?�?�?�?�?�?�O�?)OOMO;Lv�P�BPN��{��/�O 8�O�O�O_�O&__ J_5_n_Y_k_�_�_�_ �_�_�_o�Oy�Co�� LoNo`o�o�o�o�o�o �o�o8&\J�jw  2o�� ���� �2�D�V�d����������Џp�o��
 � �]OS�e�w������� ��џ�����+�{B�4���{J��$�MSKCFMAP�  -��� wvD�E� � ]�ONREL  qEt�jp]�EXCFENB��q
r�����FNCƯ���JOGOVLI�M��d����d]�K�EY����_�PAN��-�)�]�R�UN��]�S?FSPDTY�@Ȧ<����SIGN�����T1MOT����]�_CE_GRP� 1�-�t�\ ��	��-�?ϗOc�� sϙ�PϽ�t϶��Ϫ� �)��M��q߃�j� ��^߱��������� 7���[��P��H���l�]�QZ_EDI�T��n���TCOM_CFG 1�j����)�;�
��_/ARC_âqE�UAP_CPL_��դNOCHECK� ?j�  pE�����������  2DVhz�������NO_WA�IT_L����װN�UM_RSPAC�Eg���=�7A�$?ODRDSP^��ѨOFFSET_�CAR����tDI�S�rPEN_FILE���=���S�PTION_IO�#�5��M_PRGw %#%$*/�".�WORK %����hpG@S%� �mDC���m ��m!	 ����m!<����TR�G_DSBL  �-���z��/��ORIENTTO�����C���s�A �rUT_SIM_ED�q�D�TVX?LCT �#B�|@-5_PEXE�g6RATs0	�ѥx�|k2yUP �<>
%�.���?�?�?O�I�$PARAM�2೏����&3	 d��VOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�� ��_�_o#o5oGoYoko}o�o��<�_�o�o �o�o&8J\ n��^"�o�����P�
��.�@�R� d�v���������Џ� �����N�`�r� ��������̟ޟ�� �&�8�J�\�+�=��� ����ȯگ����"� 4�F�X�j�|������������߿�3���!��D�R�ĽĽ���p�� �ǰ� �ϸ��������.�DO ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }�������_���� ��1�C�U�g�y��� ���o��������	 -?Qcu���# ����x�	- ?Qcu���� ���//)/�M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? </�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�Ol�ο��O4�_ (�_P_^��O�ϛ_� 0���_�_�_oo2o H�aoso�o�o�o�o�o �o�o'9K] o�������Vo ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� �����x?ޟ�-� ?�Q�c�u��������� ϯ����)���
� _�q���������˿ݿ ���%�7�I�[�m� <�N��ϵ��������� �!�3�E�W�i�{ߍ� �߱ߤ_���O��_F_ ,�:_P�^_�߂_��_ <o����������"� Hoa�s����������� ����'9K] o������� �#5GYk} ��������/ /1/C/U/g/y/�/�/ ���̟�/�/��?-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;O
? _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _NO�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o~�����F� ,:�$bp��o�� 0�B��������D� �$PARA�M_GROUP �1�gX���L��`8� � ���q�� @D7�  ��?�����1?�p���qC>������t�  ;�	�l��	 �����Xð΀π���^� �,X ����pH��H����H�33H���H�WH-����|�#�o�oi��~�qB�  B���������������s��4  �p�����ô�����������ȟ�s�����l{uÕq������r,�2���G��wρ,[��|�|��p��?�  Д������u	'� �� ТI� ��  �����=���������@��"����F�����0��[�i���������Z��CݐB���a���B��б��Ŀֿ�   ��C9>���� :�}
<�H�wB��L�+�XŎ�� 3�tŕqDz������Ϧ�����pȯڨ�!�  �,��:=˅�!D� ?�ff{R�d��Ϗ ���ߪ���8������ڰ�D�����(����P�!�A������f�?333}���;���;QaT;�\��;��;�	�<$D4�Lq��A0s봂���?fN�q���?3�?y&����A���@�,����©� ���ɤ����#���� ��X�C�|�g������� ��������0T ?x����q�m�E�  E;��E@ Eꃂg <N9r]�� ����s�/o�./ ��a/��/��/�/��/�/�哠�?��|�3�M�A��/=?(?�a?L?�?p9A+�A� �4���!�?;�y?�?u7xo�Ϗq<?��O�OKO6OaI��3��mk^OC����`󲈣OJ(%D�%@$A�A@�I�`MD/��CG33Ck��B�1B-v��=���̞�E��ីW
Ͻu�OjC²�B����0X��Blz��X���(^�
=Õ���ö�=BU(�������E@K���JD��LU�W�H�� I%�K�A	�aLLU�L =�L]���HP� H�R���_�PTF�L%��J�
`H���H���A�� `OoL_�_7o"o[oFo ojo�o�o�o�o�o�o �o!E0iTf �������� �A�,�e�P���t��� ��я��Ώ��+�� O�:�s�^�������͟ ���ܟ� �9�$�6� o�Z���~�����ۯƯ�����5� �G�><;�A� C��3����Ć�����C�V�������޿����O�:�s�^�=(d��`��{�4������dų$rcx�Ϯ�^�3-NQ�Ϝ����v��߰�v3�g� ��2�!�;�%D93ҵ�L�Lٌ�zߠ�ߞ������5Pl�P�A"//��;�e�P��t�)�����D��������@8�0t���S�>�w�b����B�/��������9`��8&HO�H�Z  �e 3�t6�����  2 E\~C��E�`/����B���2�0C��@�0��@�?z���Q�r0 F�� G�� D	�C CE�� F��@/!/3/E/W/��?��Tp!��������r��4K
 ^/ �/�/�/�/	??-??? Q?c?u?�?�?�?���2{����uD�Y�4ӀK�&��1 @�DE�1?vPA � `?m!vT��5��2L;�	lB�}��RKLC@iK��F����2O�?�O����O�L��$H�O�O� $__H_3_l_W]E`@��_�W��_!��A���_�Xa_o]U+UU<oo=���Tofk� cv`�0�o�hb&f��o�m�2�	�o}^u0  '��vo2�]_V��B�OyAxB8U��| .�u4C�F�B�
��C�.�,b6�m�{�  �6�:�"�!� ��B>���ÏU� �����=�+� �2�>ua�0A4�y�k���I�>L~a�T=�A@�Ϻ���ۏi%	A�3|B�p?fff?.?&�9�*�6�B	� D4�Ed�H���HD �����ܯǯ ��$� �H�Z�E�~���g��� ��ؿO�q�s�ѿ2�Ϳ V�A�z�eϞωϛ��� ��������@�+��_ s�9ߚ��������U� ��*�<�۟Q�c���@���������T��iX���;�&� ϕ�o%���q������� ������(L7 p�m����� ��H3lW �{�����/ �2//V/A/z/e/w/ �/�/�/�/�/�/?? @?R?=?v?a?�?�?�? �?�?�?�?OO<O'O `OKO�OoO�O�O�O�O �O_�O&__J_5_G_ �_k_�_�_�_�_�_�_ o"ooFo1ojoUo�o yo�o�o�o�o�o�o 0T?x�u����w(�q������&��J�8� n�\�~�����ȏ���@ڏ���4�"�]�P̒	Pf���b�����x ��ş���ԟ���1� �U�@�R���v����� ӯ������`�*���3� 5�G�}�k�����ſ�� �׿����C�1�g�u�  2�ϭϿ� ��������+�=�K���o߁ߓߥ߷���8�����
 ���� D�:�L�^�p���� �������� ��b�����{J�_��+�[�H� @D��  \�?�b� �G `?��h���C]��\�X��� ;�	lh�c�}�����l�<����F�������+����.�Є� N	�߄o��� �]�����]�Y�.�@N�r��+UUwz=��ʹ�`�X���a&f/-N�[�:/~�u0  '`/ n(a�/��/�u���/�(B �/> c@� 45�!ECw� �/[?�/?j?�?�?�q�0�?�7  Ȗ2�:�S��!%h�p�<O#O�? .��YOkK�18�0�O�J> �I�p�:�?�O�/)�c>L�Sĝ0A��O DO�O<O�3h�N�h�10?fff?40?&nP�?�_�4u�iQu� �9d��_b��_SV��_ oo<o'o`oKo�ooo �o�o�o�o�o�o�o 8�_�_�_1�-� ������4�� X�C�|�g�����%ӏ ����U�yB���f� x�����;_��ß]���`���>�)�A0A�f��n�w�6��� ��/U7/���ѯ
��� �@�+�d�O���s��� ��п�Ϳ��*�� N�9�r�]�oϨϓ��� ���������8�J�5� n�Yߒ�}߶ߡ����� �����4��X�C�|� g������������ �	�B�-�?�x�c��� ���������� >)bM�q�� ����(L 7p�m���� ��/�/H/3/l/ W/�/{/�/�/�/�/�/�?�/2?7($1���T?f;P?�?t?�? �?�?�?�?�?�?(OO�LO:OpO^O�O�L��P,RP�N Q¤%?�O I8�O%__I_4_m_X_ �_|_�_�_�_�_�_o �_3ooWo�O���o� �o�o�o�o�o�o% I7Ym����w  2Ro�� �1�C�U�g�y��������Ϗ����p)�HoM�[�
 [� ;��O������П��� ��*�<�N�`�r��B�{���{J��������B�� @D��  ��?�£ �� `?>�Ȣ>�C𽤼��F� ;�	9lȢ�A}���x̠)�E�F����6���A��|���E� 䨮�i�G��Ͽ�� ,�ͽ� �Q�_ǽ��v��РϮ�!�����+UU����=����&���6и�@�N���&fd�vݮ��y���=�u0  ' �����������բ�a�9��B W��� @����EC �A���������������-�;�  �"��:o��qU��uȢ���q���� �@������8������>5ѩ�С��9�+S�Ɖ�>L>ѳt��A�@D��B����Ȣ��|Ȣ��?fff?��?&� �����բ� դ��ĥ$¨D�� �xc����� �///>/P/'/t/ _/�/13�/�/�/ ??:?%?^?I?[?�? ?�?�?�?�? O�?�� 3O�?ZO�/{O�/�OO �O�O�O�O�_#_�O�V_A_z_e_�_�_Am�A��T��S�_�_ �_�Z����_Fo1ojo Uogo�o�o�o�o�o�o �o0B-fQ� u������� ,��P�;�t�_����� ��Ώ���ݏ��:� %�7�p�[�������� ܟǟ ����6�!�Z� E�~�i�������دï ��� ��D�/�h�z� e�����¿���ѿ
� ���@�+�d�Oψ�s� �ϗ����������*� �N�9�r�]�oߨߓ� �߷��������8�J�5�n�Y��}�(�������������� 
���.��>�@�R��� v�������������e%P�P&=A"d�� V��[�p��� ��� K6 oZ�~�^ O� DH��/=/+/a/O/ �/s/�/�/�/�/�/?8�/'?7  2�[? m??�?�?�?�?�?�?�?JJ?/OAOSOeO�wO�O��O�J
  �O�G�O__0_B_ T_f_x_�_�_�_�_�_�"�O��{J���$PARAM_M�ENU ?�U��  �DEFPUL�SE�[	WAI�TTMOUT/k�RCVBo S�HELL_WRK�.$CUR_ST�YL-`nlOP3TA9a�oTB�o�b�CioR_DECSN:`�l�o�o1 ,>Pyt������	�aSSR�EL_ID  ��E1��USE_PROG %jq%�j��CCRF`�*�1c}�_HOSoT !j!����w�T7 ��ۃ�����݃�v�_TIM�EDb*���`GD�EBUG(�k�G�INP_FLMS�K@�o�TR~� �q�PGA�� _�f�I ���CH}��  q�TYPE
l@��4�]� X�j�|�������į� ����5�0�B�T�}� x�����ſ��ҿ�� ��,�U�P�b�tϝ���Ϫϼ���q�WOR�D ?		�FOLG-c	U��	MAKRO�+�SUCHL�C�2�S7T�TRACECTL 1��U�a
 �@�� ��@  {�2�ߗߩ�S�_DT Q��U���o�D � 	W� ����Г��U��ԕ�Ԗ�ԗ��U��ԙ�Ԛ�ԛ��U��ԝ�Ԟ�ԟ��U��ԡ�Ԣ�ԣ��U��ԥ�Ԧ�ԧ��U��ԩ�Ԫ�ԫ��U��ԭ�Ԯ�ԯ��U��Ա�Բ�Գ��U��Ե�Զ�Է��U��Թ�Ժ�Ի��U��Խ�Ծ�Կ��U������������U������������U������������U������������U������������U������������U������������U������������U������������U������������U������������/� ��s�B���1��P�� z������� �� ��	�
��
���� �� "� *� 2�D@dcސ� ��������J�����g%������������������G� �*���5����' ��' �' �' �����V��W��X��Y���Z��[��\��]���^��_��`��a���b��c��d��e���f��g��h��i���j��k��l��m���n��o��p��q���r��s��t��u���v��w��x��y���z��{��|��}���~���Ԁ�ԁ��Ԃ�ԃ�Ԅ�ԅ��Ԇ�Ԉ�ԉ�Ԋ��ԋ�Ԍ�ԍ�Ԏ*�ԏ�Ԑ�ԑ�����1� ��P�+H��9OKO]OoOK�uLܕOwJ�uL�!�J�M�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_vK�o'o 9oKh��YokoMo�o�o �o�o�o�o�o1 CUgy���� sO��	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ�� �%�7�I�6B'Io��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ������������ �%�7�I�[�m���� ������������! 3EWi{�{ek� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o ��o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� ��o=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?1�?�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y�����s?��ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ������������' 9K]o���� ����#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o��1oWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ����	��-�?�Q�c�u���$PGTRACE�LEN  v� � ���A`ȋ�_UP _�����������y����_CFG7 �����Aa������ĝ�����������DEF�SPD ���l@a��Ћ�IN��?TRL ������8��V�PE_CO�NFI�����������#�L�ID�á����G�RP 1���� �v�C8����VAaA��
=G� G��L�F�( A��  D	�����d��)�9��� 	 ����S�G ´��n��B�� ������������wB<h���G�Y�C� <,1 ~�^���Z��������� ��v� 9��IoZ��z����
 �C����p�@6�QA.6p�AaH��SH�� ��r���A�,eP�>V�>W�z�v����/^�!��
V�7.10beta�%  @��@_\)@0ϣ�C9A`C C{�Z!B���B!/D�  j"0�g!����� Df�� R!�B� �"C�> �� �!��� ;��B���B33B7� (�� �!B ffB�!��A�ff���˚¸��*=3���/?��C�&�8�ѩ�� [?�?j?�?�?�?�? �?�?�?!OOEO0OiO TOyO�O�O�O�O�O�O _�O/__,_e_P_�_ ܳ �_�_n_�_�_�_ oo=o(oaoLo�opo �o�o�o�o�o�./T#F@ >y:}N`|~ ?�&�� ����/�??/?A? J��on���k�����ȏ ���׏����F�1� j�U���y�����֟� ӟ���0��T�?�x� ���_����o��ϯ� �,��)�b�M���q� ����ο����1 c=�O�y���ϸ� �����	��-�?�H� �l�Wߐ�{ߍ��߱� �������2��V�h� S��w�������� ����.��R�=�v��� ����[��������� *N9r�o� �����/�a� ;Mn�ϒ������$PLID_K�NOW_M  >:%�>!�?SV �������� ��)/;/M/�q/\/n/�/�� �M_G�RP 1��� l�C9�"�g� �&�$ }0=H��@�("1 *5&?8<���	7�+a? ???�?S?e?�?�?�? 	O�?�?9O�?OuO+DV�MR�#��-T�Ί�  �"�Cf ���O�N_�O���O >___$_�_H_�_�_�~_�_�_�%ST�!1W 1��"`� �0Vacia�rC��;>�A@��A����H>y�H��hA
C/La�rguero7f����p�@Q�D�A%JvOb����H�c�Llen1lq`���p@6�QA.�6pOb��SH���V���F�o   �o�o�o�o2'h K]o�����"g2o)`� �C� �8�J�x�n�����ӏ ��ȏڏ����"�c� F�X�j����������k3�(��̟-�n� Q�c������������� ��4��)�;�M����q���Ŀ������c4 �'��˿,�m�P�b� �φϘϪϼ������� 3��(�:�Lߍ�p߂ߠ�ߦ߸���c5��&���<)�n6 �%�7�I�c7b�t����c8��������~cMAD  �$�"c  dPARNUM  ���"��7�T_S+CHN� \�
��o�8�����UPDo�����!b_CMPa_� Q���'��S_ER_CHK6���cO3�ERS�@��"_M�OP���_��R�ES_G`�� �?aC�|�%#ߛH�|������oaC�8�(B�}vH��j4�� �`D�K�HB�oH�1�T� U  NOTMqv���� ���%/XI��� 1//�/y/�/�/�/�/ �/?�/(??L???Q? p?6/��Q/�?u?�? �?	O�?-O O2OcOVO �OzO�O�O�O�O�?� ��?�O�OD_7_h_[_ �__�_�_�_�_�_
o��_o.o�O��\ _Qo�a�no�o�o� ��o�o�o����o<�V 1���������^�`��^��]����]���THR_GINR� S��d��d�vMASS� �Z�wMN��sMO�N_QUEUE ��š��ȡ��%MJ� 2��y���4A�  @���Bʡ��c*	�N- UqN�v_�m�ENDo����EcXE������BE��|y�j�OPTIOv���m�PROGRAoM %�z%l��J3�k�TASK_�IP�ߎOCFG ����󔟛�OD�ATA�1�}��@  ��? 2 �ޟ�`��&�0�ڑ F� X�j�|�����C�����pѯ���� �� ڟ*�<�N�`�4����� ����̿�����&� 8��p�nπϒϤ�x� ����������4�F� X�j�|�PϠ߲����� �߼���0�B�T�(��x������s�IN�FO���}�� �c
��.�@�R�d� v��������������� *<N`r��5I���� =is�~��DIT �}��@mU��C!OWER�FL��rs��RGA�DJ �}�A�  '?��3�q�m�x��U��?C�ѐ <@	�����%qq����I�J��U˒��\9fqrbb�A<t�t$&�* /" **: ""��/'#UL"G%#��!Q)Q��� q/sE/W/i/{/�/�/ �/�/�//?�/??�? �?S?e?w?�?�?�?�? �?�?�?OO+OUOOO aOsO�O�O�O�O�O�O �O__'_9_K_]_�_ �_�_�_�_$o�_�_�_ oko5oGoYo�o�o�o �o�o �o�o�o; 1CUg���� ����	��-�?��Q�c�u������ 	 ��,��P�;�	)u�# A���=�Ɵ���
/ /�@/ʏ܏q� ��� L�^�˯��������� ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�Dϱ�h�z� �Ϟ����������N� �.�@߭�d�v߈ߚ� ����������*� <�N�`�r����� ��������&�8�J� \�n������������� G��"4�Xj |����
C. l�v<�8�؟� ��� �2����� �>/P/b/t/�/�/�/ �/�/;?�/??(?~? L?^?p?�?�?�?�?�? 7O�? OO$ONOHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_o�_�_�_
o wo.o@oRodo�o�o�o �o�o�o�os* <N`����� �����&�8�J� \�n��������#�� G�^h����R���ş �� /*/�6/��ҏ g�����B�T�~�x��� ������ү����� ,�>�P�b�t������� ��ο�M���(�:� ��^�pςϔ��ϸ��� ��I� ��$�6ߣ�Z� l�~ߐߺߴ������� ��� �2�D�V�h�z� ������������
� ���@�R�d�v����� ������&��� <N`r����  9Kb�l���.����$PRGN�S_PREF }���� �� 
�IORI�TY  ݔ�����MPDSPON  ݖ0���#UT&��5&ODUCT_IOD �"���OGGRP_T�GL$m&V&TOE�NT 1�i*�(�!AF_INE�E �/�!tc�p�/�!ud��/�!icm�!?�Z"XY_C�FG ��+ ��)� #��?�?� ��?�?�5�?�? �?!OOOWO>O{ObO��O�O�O�O�O�O_*4Y#t3�� %�O_�a_�>�%��B#�/�:_�_��-%��X�A���,  ���_
oo.o)(T����0"��PORT_NUM�#� %�_CARTREP& |{<�SKSTAE'� �jSAVE ��i*	260_0H613���!�_'3?K !	ox����ݓ�e������
��|JU��e_�  1���+ p �*�j���#��������a_CONFIw0�Zg#�]�U�ޔy��0��}�ȃPt22�֋���[��`C�U��$�q�2�։��a����:�8��o�>�\?L���?
XH�+���?�!?���?:��>�;��C��OCe��OEn����q��UZ���������Ŕe�͔�Օٕ?����V�p�� �+�����y��� i�����_������_� �U]��A���Q�w�� ۯ�����#����Y� �=�˿)�sυ�׿� ��������U���9� Kߝϯρߓ��Ϸ��� �������c߭�G�Y� ��}���ߛ����)� s�����C�U���y������k2S_MOT�I$ 2�֋
� ?���_��);M�`�5����x����Z +=Oas�� �����y��#� &/./@/R/d/v/�/ �/�/�/�/�/�/:� /7?I?[?m??�?�? �?�?�?�?�?O
?? EOWOiO{O�O�O�O�O �O�O�O__/_*O<O e_w_�_�_�_�_�_�_ �_oo+o=o8_J_Jo �o�o�o�o�o�o�o '9K]Xojo� �������#� 5�G�Y�k�fx��� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u������������� ��)�;�M�_�q��� ��������Ư��� %�7�I�[�m�ϑϣ� ������Կ��!�3� E�W�i�{ߍߟ߱��� ���������/�A�S� e�w��������� �����=�O�a�s� �������������� �"�"]o�� ������# 50Bk}��� ����//1/C/ >Pb�/�/�/�/�/ �/�/	??-???Q?c? ^/p/�?�?�?�?�?�? OO)O;OMO_OqOl? ~?�?�O�O�O�O__ %_7_I_[_m__�_�O �O�_�_�_�_o!o3o EoWoio{o�o�o�o�Q�Q�Q�e�i%�f�o�g�4�o �A���m�c�S�e  88R�Q8_�|��� �_ �_�	��-�?�Q�c� u���������Ϗ�_� ��)�;�M�_�q��� ������˟ݟ���� %�7�I�[�m������ ��ǯٯ�����
�
� E�W�i�{�������ÿ տ������*�S� e�wωϛϭϿ����� ����+�&�8�J�s� �ߗߩ߻�������� �'�9�K�F�X߁�� ������������#� 5�G�Y�T�f�x���� ��������1C Ugyt������ ��	-?Qc u������� //)/;/M/_/q/�/ �/�/���/�/?? %?7?I?[?m??�?�? �?�?�/�/�?O!O3O EOWOiO{O�O�O�O�O �O�?�?�O_/_A_S_ e_w_�_�_�_�_�_�_ �_�O_+o=oOoaoso �o�o�o�o�o�o�o �_o"oK]o�� �������#� 0Y�k�}������� ŏ׏�����1�,� >�P�y���������ӟ ���	��-�?�Q�L� ^���������ϯ�� ��)�;�M�_�q�l� ~�����˿ݿ��� %�7�I�[�m��z��� �����������!�3� E�W�i�{ߍߟߪì��������%������'���������Ӡ���  (�B���8O����� �Ϯ����� ��/�A�S�e�w��� ������������ +=Oas��� �������'9 K]o����� �����5/G/Y/ k/}/�/�/�/�/�/�/ �/?//C?U?g?y? �?�?�?�?�?�?�?	O O?(?:?cOuO�O�O �O�O�O�O�O__)_ ;_6OHOq_�_�_�_�_ �_�_�_oo%o7oIo D_V_h_�o�o�o�o�o �o�o!3EWi dovo������ ��/�A�S�e�w��� ����я����� +�=�O�a�s������� ��͟ߟ���'�9� K�]�o����������� ğ����#�5�G�Y� k�}�������ſ��ү ҿ��1�C�U�g�y� �ϝϯ��������� �-�?�Q�c�u߇ߙ� �߽��������� �� ;�M�_�q����� ��������� �I� [�m������������ ����!�.�@�i {������� /A<Nw� ������// +/=/O/a/\n�/�/ �/�/�/�/??'?9? K?]?o?j/|/�?�?�? �?�?�?O#O5OGOYO kO}O�O�3�1�1�E�I%�F�O�H�O�O�Ox�E�3�E  _2_�18?_u_�_>�_� �?�? �_�_�_oo1oCoUo goyo�o�o�o�?�_�o �o	-?Qcu ������o�o� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ�����
�3�E� W�i�{�������ïկ ������*�S�e� w���������ѿ��� ��+�&�8�a�sυ� �ϩϻ��������� '�9�4�F�Xρߓߥ� �����������#�5� G�Y�T�fߏ����� ��������1�C�U� g�y�t��������� ��	-?Qcu ��������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ ���/�/?!?3?E? W?i?{?�?�?�?�?�? �/�/OO/OAOSOeO wO�O�O�O�O�O�O�? �?O+_=_O_a_s_�_ �_�_�_�_�_�_o�O _9oKo]ooo�o�o�o �o�o�o�o�ooo 0oYk}���� �����1�,> g�y���������ӏ� ��	��-�?�Q�L�^� ��������ϟ��� �)�;�M�_�Z�l��� ����˯ݯ���%� 7�I�[�m��������Ę���%����Ƕ2 y���� �Ĥ�x������  �"ς�8/�e�w�>��� |��� ���������!�3�E� W�i�{ߍߟ�r����� ������/�A�S�e� w���������� ��+�=�O�a�s��� �������������� '9K]o��� ��������#5 GYk}���� ����C/U/ g/y/�/�/�/�/�/�/ �/	??/(/Q?c?u? �?�?�?�?�?�?�?O O)O$?6?H?qO�O�O �O�O�O�O�O__%_ 7_I_DOVO_�_�_�_ �_�_�_�_o!o3oEo Woiod_v_�o�o�o�o �o�o/ASe wro�o����� ��+�=�O�a�s��� ����͏ߏ��� '�9�K�]�o������� ����������#�5� G�Y�k�}�������ů ��ҟ����1�C�U� g�y���������ӿί ���-�?�Q�c�u� �ϙϫϽ��������  �)�;�M�_�q߃ߕ� �߹�����������  �I�[�m����� ���������!��.� W�i�{����������� ����/A<�N� w������� +=OJ\� ������// '/9/K/]/o/z|rD�%�)%�&�/�(�/�/ EAL�-�#p�%  �/?r�8?U?g?y?� l~�?�? �?�?�?O#O5OGOYO kO}O�Ob�?�O�O�O �O__1_C_U_g_y_ �_�_�_�O�O�_�_	o o-o?oQocouo�o�o �o�o�_�_�o) ;M_q���� ���o�o�%�7�I� [�m��������Ǐُ ���
�3�E�W�i� {�������ß՟��� ���A�S�e�w��� ������ѯ����� �&�8�a�s������� ��Ϳ߿���'�9� 4�F�oρϓϥϷ��� �������#�5�G�Y� T�fϏߡ߳������� ����1�C�U�g�b� tߝ����������	� �-�?�Q�c�u����� ���������) ;M_q������ ���%7I [m����� ��/!/3/E/W/i/ {/�/�/�/�/��� ??/?A?S?e?w?�? �?�?�?�?�?�/�/O +O=OOOaOsO�O�O�O �O�O�O�O�?�?O9_ K_]_o_�_�_�_�_�_ �_�_�_o__GoYo ko}o�o�o�o�o�o�o �o1,o>ogy �������	� �-�?�:Lu����� ����Ϗ����)� ;�M�_�j�l�b�x���q%s�����'"���͟o�����`��� � ��b�8��E�W�i�� \�n�����˯ݯ� ��%�7�I�[�m�� R�����ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭ߨ� �Ϻ�����+�=�O� a�s��������� ����'�9�K�]�o� ���������������� ��#5GYk}� �������� 1CUgy��� ����	/( Q/c/u/�/�/�/�/�/ �/�/??)?$/6/_? q?�?�?�?�?�?�?�? OO%O7OIOD?V?O �O�O�O�O�O�O�O_ !_3_E_W_ROdO�_�_ �_�_�_�_�_oo/o AoSoeowor_�_�o�o �o�o�o+=O as��o�o��� ���'�9�K�]�o� ��������ۏ��� �#�5�G�Y�k�}��� ��������ҏ���� 1�C�U�g�y������� ��ӯΟ��	��-�?� Q�c�u���������Ͽ �ܯ� �)�;�M�_� qσϕϧϹ������� ����7�I�[�m�� �ߣߵ���������� !��.�W�i�{��� ������������/� *�<�e�w��������� ������+=O Z�\�R�ht	%c�Η�[��� ���ttP�t � ��R�8��5GY� L�^������ �//'/9/K/]/o/ B�|�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �/�/�?�?�?�?OO 1OCOUOgOyO�O�O�? �?�O�O�O	__-_?_ Q_c_u_�_�_�_�_�O �O�_oo)o;oMo_o qo�o�o�o�o�o�_�_ �_%7I[m �������o�o !�3�E�W�i�{����� ��ÏՏ������ A�S�e�w��������� џ������&�O� a�s���������ͯ߯ ���'�9�4�F�o� ��������ɿۿ��� �#�5�G�B�T�}Ϗ� �ϳ����������� 1�C�U�g�b�tϝ߯� ��������	��-�?� Q�c�u�p߂߂���� ������)�;�M�_� q�������������� %7I[m ���������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/���?+?=?O? a?s?�?�?�?�?�?�? �?�/�/'O9OKO]OoO �O�O�O�O�O�O�O�O _OOG_Y_k_}_�_ �_�_�_�_�_�_oo _,_Uogoyo�o�o�o �o�o�o�o	-? JcLaBaXudy%Sv}·vU
�t� �� d}ds@cdu � ��Ba8��%�7�I�� <oNo��������Ϗ ����)�;�M�_� 2ol�������˟ݟ� ��%�7�I�[�m�� z�����ǯٯ���� !�3�E�W�i�{����� ����տ�����/� A�S�e�wωϛϭϨ� ��������+�=�O� a�s߅ߗߩ߻߶��� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ��������������� 1CUgy��� ����	? Qcu����� ��//)/$6_/ q/�/�/�/�/�/�/�/ ??%?7?2/D/m?? �?�?�?�?�?�?�?O !O3OEOWOR?d?�O�O �O�O�O�O�O__/_ A_S_e_`OrOr_�_�_ �_�_�_oo+o=oOo aoso�o�_�_�o�o�o �o'9K]o ���o�o�o��� �#�5�G�Y�k�}��� ����������� 1�C�U�g�y������� ����Ώ��	��-�?� Q�c�u���������ϯ �ܟ��)�;�M�_� q���������˿ݿ� ����7�I�[�m�� �ϣϵ���������� 
��E�W�i�{ߍߟ� ������������/� :�<�2�H�T�%C�m�z�d��P�V�0�T� � ����2�8����'�9�� ,�>�w������� ��������+= O"�\������ ��'9K] oj|����� �/#/5/G/Y/k/}/ x��/�/�/�/�/? ?1?C?U?g?y?�?�? �/�/�?�?�?	OO-O ?OQOcOuO�O�O�O�? �?�?�O__)_;_M_ __q_�_�_�_�_�_�O �Ooo%o7oIo[omo o�o�o�o�o�o�_�_ �_!3EWi{� �������o /�A�S�e�w������� ��я������&� O�a�s���������͟ ߟ���'�"�4�]� o���������ɯۯ� ���#�5�G�B�T�}� ������ſ׿���� �1�C�U�P�b�bϝ� ����������	��-� ?�Q�c�u�pςϫ߽� ��������)�;�M� _�q��~ߐߢ����� ����%�7�I�[�m� �������������� !3EWi{� ��������� /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ �/�/��'?9?K?]? o?�?�?�?�?�?�?�? �?�/?5OGOYOkO}O �O�O�O�O�O�O�O_�_���$PUR�GE_ENBL � ,A-A��-A4PWF<PDOG  DT,BOQ TRS_I]TgQKUTQ�RUP_DELAY �"A"AKU,B��R_HOT %��UiR%+B�_�]�SNORMAL�XKR�_<!o�WSEMI o&o�eopQQSKIP_�GRP 1ĞU�MQ x 	 ho�o�o�o�o�o�i �U'wGYk1 �}������ �1�C�U��e���y� ����ӏ������-� ?�Q��u�c������� ��͟���)�;��U�$RBTIF^T��ZY�CVTMOU�T^V�U�Y�D�CR�cƈi ���aEVQ�E��2E�npD�&�DFoFC��3[�m�R�,��ֶ�&���b��ĆB�×�	�o� �;��;Qa�T;\��;���;�	�<$�D�/@�j�{� {�����ſ׿��� ��1�C�U�g����� vϯϚϿ�����	�L� -�?߂�c�u߇ߙ߫� ����������)�;� ��_�J��n���� �� ���V�7�I�[� m�������������� ������3WB{ f������*� /ASew�����,kRDIO�_TYPE  �[��REFP�OS1 1Ǟ[
' xSoY)�}/ ��/�-L/^/�/�/�/ ?�/A?�/e? ?b?�? 6?�?Z?�?~?OO�? �? OaOLO�O O�ODO �OhO�O_�O'_�OK_ �Oo_�__._h_�_�_ �_�_o�_5o�_2oko o�o*o�oNo�o�o/%/2 1�;+J/�o �oL�opvo�/� ������6��xZ�l�-'3 1� 
��V�ԏ������ ��@�ۏ=�v����5�ྟY��p�0$4 1ʍ�����۟Y�D�}� ����<�ů`�¯��������C�ޯg���0$5 1���&�`�޿ ɿ��&���J��G� ��Ϥ�?���c���z�^0$6 1�;+�������`��τ��3!7 1��.�@�z��������S8 1� ��������x��/��SMASK 1��� H ������XN)O���4�D�/!?MOTE  �M�_CFG �[��D�."PL_RAN�GW�+!_���OW_ER �;%���g�."SM_DRY�PRG %;*%�X� ��TART ����
UME_�PRO����j,$_�EXEC_ENB�  �c�GSP1DC � �e���GTDB��
RM\��MT_��T���Y��OBOT_I/SOLC�����x'NAME �;*KJLT�VL411550wR01x2 0#�_ORD_NUM� ?��
!H613 ��_895 ܶ\��P+!�  ������� 8�/ PC_TIME�OUT�� x/ S7232t�1�;%�� LTEA�CH PENDA�N�p�G�I�n�W��Maint�enance C�onso�C�R,"�b/��	UnbenutztY*�/X/�/��/�/�/�/�b"NPqO �K����SCH_LF ����	�1T;MA�VAIL��5���c�SPACE1 {2��
 K?@HHG�v�F�������4L8�?� L;WOL?;O�O�O�O�O �G�?OO%O�OIOkO ]_~_A_�O�_�Y�#� �]�O__%_�_I_k_ ]o~oAo�_�o�o�o�O �_o!o�oEogoYz =�����o�o /�Suw9��� ����������+� ُO�q�c��������� ��ߏ���'�՟K� m�_���3�������˯ ����#�ѯG�i�[� |�?�������ǿ��� ��1�C�U�WϾ�;� �Ϯυ������	�� -���Q�s�e�7߉ߪ��ߓߥ��52�?�?�� �#���G�i�x��\� ����������*�<� N�`�r�t���X����� ������&�8�J��� n����T���� ��"4F�j� ~�R���� 0B�f�z/�/ ^/��/�/�///,/ >/�/b/�/v?�?Z?�? �?�?�???(?:?L? �?p?�?�?VO�O�O�O �O OO$O6OHO�OlO �O�_�O�_�_�_�_�O _ _2_D_�_h_�_|o �oPo�_�o�o�o
oo .o@o�odo�ox�\ ������3��
� .@�d����� y�ˏ�ӏ�5�G� Y�k�}�������u�ǟ 蟿����1�C�U�g� �������q�ï��� ͯ�-�?�Q�c���� ������o����ٿ� )�;�M�_�σ����� ��{�ݿ�����%�7� I�[�	�ϡϓߴ�w� ��������!�3�E�W� i��߯߱�s����� �����/�A�S�e�� �������������� �+�=�O�a����� ��m����' 9K]����@y���/�4� '�9K]/���/ �/�/�/	?�/?#R/ d/v/�/�/�/�??�? �?O�?O<?N?`?r? �?2O�?�?�O�O�O_ _�O8OJO\OnO�O._ �O�O�__�_�_o�_ $oF_X_j_|_*o�_�_ �o�o�o�_�o Bo Tofoxo&�o�o�� �����>Pb t�4������� �ڏ�:�L�^�p��� 0���ȏ���ޟ��� ��6�H�Z�l�~�,��� ğ��ׯ�������"� D�V�h�z�(��������ӿ���	���#+52.D/V�h�z�(Ϟ� �����ϳ��&��;�#+6O�a�sυϗ�E� ���������"�C�*�X�#+7l�~ߐߢߴ� b�����	�*���?�`�G�u�#+8����� ������&G
\�}d�#+G �N5+ �:
�  �,: 5%K]o������ ��o�>d � %/7/I/<j/|/�/�/ ����*�/�+?
/ ;?M?_?q?d/�?�?�? �/�/�/�/?O7O*? [OmOO�O�?�O�O�O��?�?�?O$O6_ `� @> oU� }_�O�_�Ek_9_�_-O o�_�_�_�_loo1o So�ogo�A�a�E�c�o �o!�e�oSe �9k���������L
�_n�@��_MODE  ����S ��]�_Z���_��9�	4�]�D�CWO�RK_AD���{9�F�R  ����b���_INOTVAL��������R_OPTION�̖ ��F�TC�F� ۗ���?���7���V_DATA_GRP 2��H�DU@PJ�y�F� ����G�ʯ���ܯ�  �6�$�F�H�Z���~� ����ؿƿ����2�  �V�D�z�hϞόϮ� ���������
�@�.� d�R�tߚ߈߾߬��� �������*�`�N� ��r��������� ��&��J�8�n�\�~� �������������� 4"DjX��Be� �������q�5 #YG}k��� ����//C/1/ O/U/g/�/�/�/�/�/ �/	?�/??-?c?Q? �?u?�?�?�?�?�?O �?)OOMO;OqO_O�O �O�O�O�O�O�O__ _%_7_m_[_�__�_ �_�_�_�_�_�_3o!o WoEo{oio�o�o�o�o ��o� ��o�oA we������ ���=�+�a�O��� s�������ߏ͏�� '��3�9�K���o��� ��ɟ���۟����� G�5�k�Y���}����� ���ׯ���1��U� C�e�g�y�����ӿ�� ����	��Q�?�u� cϙχϽϫ������� ��o>�b�M�ߕ� ߹ߧ��������� �%�[�I��m��� ���������!��E� 3�i�W�y�{������� ������/e S�w����� ��+O=sa ������/ /9/'/I/K/]/�/�/ �/�/�/�/�/�/�/5?�#?Y?+��$SAF�_DO_PULS�  -��������1t0CA?N_TIME�0}���3���1R ������8�		����
�8����4�4��  ^�OO0OBOTOfO�?��O�O�O�O�O�O�G��1  B2�T�1�1dXQ Q��4}��1�� @ CVT[�0P_z_�\�1�_��WP�U�� {@B�3T i_��_�_oiT D��oAoSoeowo�o �o�o�o�o�o�o�+=OaX^?VNV{py 
�q�p��y�3�1;��o}��4p{}
�t� �Di�0��A�1�z   ��B�1�q�1�A�1�z�Y�k�}�������  ��������  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v���������@Я�����$��h_ H�Z�l�~�������ƿؿ'�>T�Q���R �7�I�[�m�ϑϣ�Žρ�0�22�@U<�}����$�6�H�Z�
��^�^ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x�������������� ,>Pbt� ��#�����`(:L�2��P+�imih��0�A�B Ѓ�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?OO*O<ONO#�� =X��*`YO�O�O�O�O �O�O__&_8_J_\_@n_�_�_�_�_�Z�B��_�V�_i���A��_/m	12�345678�r�`!B  �
/h�@��jo|o�o �o�o�o�o�o�o q�O #5GYk}�� �������1� C�T�w��������� я�����+�=�O��a�s�����V�BH ��П�����*�<� N�`�r���������̯xޯ�[�;�j�� &�8�J�\�n������� ��ȿڿ����"�4�F�]�D�_wωϛϭ� ����������+�=� O�a�s߅ߗ�Z����� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1C�gy�� �����	-�?Qcu���U g`���`�//n%(C��A�_J_   �mH2qB�gb%)
�Pdq#�?`��R2��/�/X�/�/�+pM$ZO���/0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O? �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_��_�_�_ ooG!�$�SCR_GRP �1���� t �G!� R%	 �Ra� Zbkbdd�f%f!�ek�wg�o�o�o(-��a �bD�` D��@ =qcw�k<�R-2000iB�/185L 56/7890� @u� �RJqOpC#
V?06.10 zp�hQKaq$�y�vZa��fIa�cIa3f!�ahj�a�y	�r�
���.�@�P���HшZ`�t^g�vO���v�{�D�*[E:r7���� ����BI�z0vaA�����G�9Bo�������4 dB�G��P�  ?����~�LD?�E:pVZ`�OG!�o��o1�.'"��受hB���B��ffB�33B�  ��ǐ���L ��c   q��va@��� ˟р��v�: 򟨛vaF@ F�`� %��I�4�m�X�}��� ��ǯ���n�����0��%�7�B�E�گ ��v�����ӿ��п	� ��-��Q�<�u��/�� �c�o����i
����8̅��Ѻ�� ߘg�Ο@�B�P�1234Ns`׀h���C$A?РƳ�㏛cd!%2�rG! ��������2�>�P�� Pv�(|����� Ibp`�t Z`�}�{yi��gϩo�i 7��P�����7uIndepe���nt Axes Qs	����n�f�w ��s�w3i��r��� j|����c��	 �n�'9��Z�� ~��S��/�� ����/���F/藦� t/��/��/�/�/�/ ?�/?=?(?a?P�:� p?�?�?Z��?R?O�? 'OOKO6OoOZOlO�O �O�O�O�O����#_f� ����k_}_�_.�Rٺ_\�n�~�o��L$o 7o��boto�oUo�o�o��o�o�o��S �����_��:�� ._������������� ��p�$6HZߏ ���'����o� ~������Hohퟀ� �#��G��h�
/�� ./P/R/d/���0� 1��U�@�e���v��� ��ӿ�?�?�����? Q�Ŀu�`ϙτϽϨ� ��������;�&�_� 
�_m��F_X_����@�_�_�_�_�V�_ w�o������o���� ���+�=��a�s���$6xBT��� �3��W��� ,�>�P�b�������� ��ΏSew��:� L�^����//+/�� ܟa/��/�/6��/Z� �/~� ?��įƯدZ? |/�?�/�?�?�?�?�? �?�?#OOGO6� �VO hOzO@��O8O�O�O_ �O1__A_g_R_�_v_ �_�_�_~���_L�� ��Qocouo�2�8�J�8ff��o��4/ Z�Wi8y���������$SE�L_DEFAUL�T  �����P�MI�POWERFL � 6e.�7�WF�DO#� .��R�VENT 1�����,��`L!�DUM_EIP�����j!AF�_INE"�Ə�T!'FT�������9!�>� ��e��!RPC_MAINf�H��T���x�'VIS��G������o!TP�PU���d�I�!
PM�ON_PROXYJ���e8����c����f���!RDMO_SRV⯯�gЯ�-�!RZ�I���h,�y�!
z�M�����ih�ſ!RLSgYNCƿ�8��>�!ROS��8���4 �]�!
CE>�MTCOM^ϲ��kLϩ�!	r�CONS�ϱ�l����,� ������B�g�.ߋ� R߯�v��ߚ��߾������?����RVI�CE_KL ?%��� (%SVCPRG1r���2����3�����4
����52�7���6Z�_���7�������8������9���� ��D������'���� O����w��$���� L����t����� ����?����g�� ���=���e��� �/��//���W/ ��/��-�/��U �/��}�/��w�� �����B?�?��?�? �?�?�?�?�?OO?O QO<OuO`O�O�O�O�O �O�O�O__;_&___ J_�_n_�_�_�_�_�_ o�_%ooIo4o[oo jo�o�o�o�o�o�o !E0iT�x�������M:_�DEV ����MC:���>�%�~�L  � ���i��!�OU�T�`�:�!�REC� 1�d5L�� �  �K 	 ��t" � �#ń! ����􍶃 ���
��	���J��D��
 �X�~�6� �>M�'�  �  $�>�a  �d5��涂�
�� � W  ��M���+ n7�� �O	�7�� �1�������� �Q �����:��<�����X��5�]����8�U-M�� �M�� �Q��U�2�� �;S�V-� � �D7��L��7�� �6U� e���?  H��V��
�����	�
 �G �U5�|�c���V4��M�� �jٯ
g�E7��q� �|�7���������g�W��.��r����Vsa�� �`�	�5��H� ��p��̑m��E)��{V9��� ��7��7������<��x��
�������y�o�Q��D	��P�M�Đԡ$� 51!���K��� �C�Z �տ�� �7�e�7�W7�m 1ϫ m��M��
�^�  �����$� ��������*K�$M� ����#Y�k��u�߫���M�bM����W�����!�E �Z̐]� ���r-�f �IM���*��D� ���)�7��2��M��ZT����\��&�A ��*M�M ����p�ߛҦ̠&M�� ���	����V�߳�ȑJ����F��@����VǡF]��X���� (����S���7�d ��=���!�� j7��� UL7��7��7��	�� T�HM�77�,��� � ��v�@V�� ������}`T��  �1�� �̡K4��� +�7�� �D���7��l��]���!�\ �?�I7����
�V��L��H������M��� ��
�޵���� p� ��I�A F7�h�Z�7��7�� �/����$��v��*����'� �i	U#!����iw��� ��f �����"7���=��� �� �����]��_���m�'=H�#D�?�(� ����P�� T�)K4������ ����x�3� �8f��۱ E 	���*�� 7�ù�u�����K4D ����E/'9s� (���ᐞ�鑹
!{�a��e��,�  "�/7���,��� ����/��4����� ��)��+��Q�	ᐷ����N� }��!/ ���8/r/_�B �3 	��?/�/��q� ��KRᐡᐧ���z�`��!+�4t��?��K�4W�Ĝ?�#��?���� @�[ᐓ���A�eAy?��O���O���� Ī��� �v��w7�� ��%�sOI�[�m�� ���]�o߁ߓߥ��_ ��������ُ�o%� �o*'`S�MmMi ������� ��!�3�i�W���{� ��Ï���Տ���� �/�e�G�u������� ���џ����=�+� a�O�q����������� �߯��9�'�]�o� Q������������ۿ �#��G�5�k�YϏ� }ϟ��ϧ�������� �C�1�g�y�[ߝߋ� �߯��������q� Q�?�u�c������ ��������)��M�;� q���e����������� ����%5[I m������� !1WE{]o ������/// /S/A/c/e/w/�/�/ �/�/�/?�/+??O? =?_?�?g?�?�?�?�? �?O�?'O9OO]OKO �OoO�O�O�O�OI_ E&__J_5_G_�_3� �O�_�_�_�_�_�_o 1ooUoCoeo�oyo�o �o�o�o�o	�o- Q?a�i��� ����)�;��_� M���q�������ݏ�� ���7�%�[�I�� ��s�����ٟǟ�� ��3��'�i�W���{� ����կ�ɯ���� �/�e�S�����}��� ���ѿ�����O�_ )�s�aϗυϻϩ��� ������%�K�9�o� ]ߓߥ߇��߷����� ���!�G�)�W�Y�k� ������������� �C�1�S�U�g���� ����������	? Q3uc���� ����)M; q_������ ��%//I/[/=// m/�/�/�/�/�/A�k_ $?g_H?3?l?W?|?�? U��/�?�?�?�?OO AOSO5OwOeO�O�O�O �O�O�O_�O+__O_ =_s_a_�_�_�_�_�_ �_o�_'ooKo]o?o �ooo�o�o�o�o�o�o �o#YG}k �������� ��U�7�e���y��� ��ӏ����	��-�� Q�?�a���u������� �ϟ��)��M�? �?K���������ݯ˯ ����7�%�G�I�[� �����ǿ���ٿ� ��3�!�C�i�Kύ�{� ���ϱ��������� A�/�e�S߉�wߙ߿� ����������=�+� a�s�U������� �������%�K�9�o� ]��������������� ��!G5kM_ ��������$SERV_RoV 1�	8��0(	\�n����!3TOP10� 1�=
 6W q�  2q��!6�E �q�6 &"$�q�. �*!��Y�PE  q���Hq�1HEL�L_CFG �p�t&�0�? �?|�/q�%RSR�/ �/�/??:?%?^?I? �?m??�?�?�?�? O��?$O5MDD<I�  �E%5OvO�OCE?Mq��O�B�@K�D\D!d�O�q��)}&HK 1�+("�O?_:_L_ ^_�_�_�_�_�_�_�_ �_oo$o6o_oZolo�~oz)OMM ���/�o|"FTOV_�ENBi$Et*OW_REG_UI�o~{"IMWAIT�b��I{OUTv�DyTIMu���WVAL,s_UNIT�c�vt%Q�LCpTRYw�t%1MB_HD�DN 2�k ( ����� >�5�G�t�k�}������̌�qON_ALI_AS ?e�iLhep���(�:�L� D��w�������X�џ �����ğ=�O�a� s���0�����ͯ߯� ���'�9�K���\��� ������b�ۿ���� #�οG�Y�k�}Ϗ�:� ���������Ϧ��1� C�U� �yߋߝ߯��� l�����	��-���Q� c�u���D������ ����)�;�M�_�
� ����������v��� %7��[m� �N�����! 3EWi��� ����////A/ �e/w/�/�/F/�/�/ �/�/?�/+?=?O?a? s??�?�?�?�?�?�? OO'O9OKO�?oO�O �O�OPO�O�O�O�O_ �O5_G_Y_k_}_(_�_ �_�_�_�_�_oo1o Co�_Toyo�o�o�oZo �o�o�o	�o?Q cu�2���� ���)�;�M��q� ��������d�ݏ����%�Ѓ�$SMO�N_DEFPRO ���N�� *SYSTEM*Ё��>�RECAL�L ?}N� ( �}׏����ԟ��� ���/�A�S� e�w�
�������ѯ� �����+�=�O�a�s� �������Ϳ߿񿄿 �'�9�K�]�o�ϓ� �Ϸ������π��#� 5�G�Y�k��Ϗߡ߳� ������|����1�C� U�g�y�������� ������-�?�Q�c� u�������������� ��);M_q ������� %7I[m �� ����~/!/3/ E/W/i/�z/�/�/�/ �/�/�/�/?/?A?S? e?w?
?�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O�O _'_9_K_]_o__�_ �_�_�_�_�_�_o#o 5oGoYoko�_�o�o�o �o�o�o|o�o1C Ugy���� ����-�?�Q�c� u��������Ϗ�� ���)�;�M�_�q�� ������˟ݟ�� %�7�I�[�m� ����� ��ǯٯ�~��!�3� E�W�i���z�����ÿ տ������/�A�S� e�w�
ϛϭϿ����� �ψ��+�=�O�a�s����$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1z� �?��%����0��� �c��G���Z?6�w���O�f����o�o������q"���֟����7�ֿ L&�g������V�����vq������������5�& �,c?>W��O��Ć��h�� ������%�����F)��6w��Z���������	�/��?��6/ �O�O&/g/��T��/"x����/�v�/b�����&? �Ϡe V?��K?�?ӄv?�?� �c�?�?�:"1 �?O֊��FO� �pP6OwO����fO�O�����O�O��1�_ ��/K/�O7_�!�&_g_YH�V_�_�c%_�_��-Q�_��_�
��?&o �cZoWo ��bFo�o�<��vo�o�G�x��o�oJ���o���u?F��l8�v ���
f��
��O� �?*��� ׶U/6���T8�f� ���V�����7��/Ə �޳�����J�E?&� ��c���W���O��� ׬5��XJ8�_� ��?�֟���_t_�G�9h6�w� מ�f����ǯ<���ׯ�ȿ�Ư�:�fE�6� ����&�g��W�V���W .��ǿ��?̶���j?�-ώЋ�l�W� �%�hFχ� ��PARAM ��{�� �	�EP���ʟ�����OFT_KB_C�FG���Չ�OP�IN_SIM  ����=�O�a������RVQSTP_DSB&��߷辪�SR �)�� � & FO�LGE011 .<����0001�������THI_CHA�NGE  �����GRPNU�M� �OP_?ON_ERR��~I�PTN )վ�C�R?ING_PR1�U����VDT+� 1y�ɢ�  	�� �����������0� B�T�f����������� ������,SP bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?k?h?z?�?�?�? �?�?�?�?
O1O.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\o�o�o �o�o�o�o�o�o�o "IFXj|�� �������0� B�T�f�x�������Տ ҏ�����,�>�P��b�t������VPRG_COUNT���|��ƒENBđ���M�4���UP�D 1���T  
����B�T�f��� ������ׯү���� �,�>�g�b�t����� ����ο�����?� :�L�^χςϔϦ��� ��������$�6�_� Z�l�~ߧߢߴ����� �����7�2�D�V�� z������������ 
��.�W�R�d�v��� ������������/ *<Nwr��� ���&O J\n����������_CTRL/_NUMГ!��!"GUN%" 2}�0��  1$ !!f%#d'o/e&��/�/�/�/ÐYS�DEBUGА1��� d�� SP_PwASSЕB?;�LOG �0��� J1�^���k$[=�c%UD1:\04.12o_MPC6? 1$(�)]?o5x82�?�2?SAV �9=�!nn- x8SV�;�TEM_TIME� 1�R+ ( w@J�"/�=�� '�^�>hF�UFsG�vO�O�@P�Ox�O�O �T1SVG YS+�ѕ'��P�ASK_OPTICONА0��ߑ'Q�_DI0�ߔTBCCFG �R+r�=�.�_`�_ ���!�_�_�_o�_5o  oYoDo}oho�o�o�o �o�o�o�o
C. @yd������	��%�6�� i�{��X�����Տ�� ���0��=P�!�G� 5�k�Y���}�����ß şן���1��U�C� y�g�������ӯ���� ��	�+�-�?�u�[� F�������˿ݿ[�� ��7�%�[�m��M� �ϑ��ϵ��������� �E�3�i�Wߍ�{߱� �����������/�� S�A�c�e�w����� �������+�=���a� O�q������������� ��'K9[] o������ �!G5kY�} �����/�1/ ��I/[/y/�/�//�/ �/�/�/�/?-???? c?Q?�?u?�?�?�?�? �?O�?)OOMO;OqO _O�O�O�O�O�O�O�O __#_%_7_m_[_�_ G/�_�_�_�_�_{_!o o1oWoEo{o�o�omo �o�o�o�o�o /eS�w��� ����+��O�=� s�a�������͏��� �_	��9�K�]�ۏ�� o�������۟���͟ #��G�5�k�Y�{�}� ��ů���ׯ���1� �A�g�U���y����� ӿ������-��Q� �i�{ϙϫϽ�;��� ������;�M�_�-� ��qߧߕ��߹����� ��%��I�7�m�[�� ������������ 3�!�C�E�W���{��� g���������A�/Qwe��� ��$TBCSG_G�RP 2���  �� 
 ?�   ���>(: t^������ ���/,//P/:/ t/�/l/�/�/�/�/�/ ?�/(?:?$?^?D?n? �?~?�?�?�?�?�?O��?6OHMA��*S�YSTEM*� V8.2306 qC�4/2x@014 A t  _F�_GF�� PARA�M_T   ��$MC_MA�X_TRQ��$^�D_MGN�CC� {AV�ISTAL�I�BRK�INOLD��FSHORTMO�_LIM	Z�M�EJ\PTPL1CU2CUU3CU4CU5CU6CUu7CU8�A h�A|��A� �__ACCEJR�W<TQ�SPATH�W�Q��S�Q_RATIO��B�S�@ 2  �	$CNT_SCwALE	ZSCL�C{IN�Q_UCA���bCAT_UM�%hYC_ID 3	*cB`_EKPGj�TPGj]PG`PAYL�OAWJ2L_U�PR_ANG�fL�W�k�a�i�a�ER_F2LSHRT�gLO�da�g)c�g)c?ACRL_Shp�gzd�BHVA` � $H�B:rF�LEX7s��@J�b�@ :$.aLENKQguTQ$DEjx�t|s�R��X�p�zSLOW_�AXIq$F1*aI�s2�x1�q�u��wMOVE_TI�Md_INERT�I%`:p	$D	�TORQUE�Q!��p��IHPACEMN��`��P�s�E^�V��p�A/�x�@�x�TCV���@��A��������@T.��@��J�A����M	�(a�>(`J_MODa�pN� R�@�gq%2�@P�^�Eo�0`$J��Xp�A�RU�F?�JK.�����KKS�VKTSVK]SJJ�0�KSJJTSJJ�]SAAKSAATSA�A
�fSAAoS�AN�1ǌ<����@�@PEw_NUQr�Vq�CFG�A � $GROUP�@�SK&cB_CON�FLIC�dB_R?EQUIRE.q�q�BU sUPDAT��v� �ELk� �ͥ��$TJ��P�JE�@CTYRa�qTN	�F˦���HAND_VB�8rVqOP�U �$]�F2�F
�TSC�OMP_SW&a ���@�F� '$$M�`�IR�C|���A��x��R��A_�}b�FDļ�MA�LA��LA�KA [Ұ�KD��LD�KD [P�PGR�Gp�ST�Gp��IZp�NXDY�`R�@ �E��ڵ�` `�g�q�g �a�g0�<Q@��p��UPKUTU]UfUoUxU�U�RVr�T r�Wt�R %�n�TP�y�ASYM�U:p�� �V�Pm�ao_SHo�g4d]��C� >oPoboto�cJ�l>P��j^�T�i
�_VI�&���Ѫ�V_UCNI�c��TS�aJ�� ������l���e��� �m�y>P1a����GtOs �T�CPPIR�A } ��ENABL�p�����$TCDE�LAY�ST��SP�EE4P  X ��I�Nڠސ��ڠGP����Q���q��@MPڢPROG9_���YPEڡ��_z�	 |�m���SE s��m���' Ǧ�WARNI��EN&���OTF�qj��3_T���MAARSuCW�\��SPDz��
 ������EA�RTBE���ET芠z���PPARGAT��FLG�u�|sUS�@E�@R&��6�%�aos6RE�AJVXTR�O;UT�A p렜��� E�̢�ID`�(d^�Uc�A� `��޵�G�Q# �PH���<��{�I�$DO�  s���z� �
�I��A��J �p0��W#�۠���q�� � T�M�ES���R���T� P��"@Pl� ��#��(�!�)T"�m�� $DUMM�Y1]Q$PS_f�pRF�pg@$�&��FLA|��2>�GLB_Tu�k�*5��b�)���8!������QSTT���SBR�PM21�_V�T$SV_�ER�`O�p3�3C�LD0p2A^����G�L��EW�A 4l��$��$Zݲ!W�3���`P�As %b� ��3U�5 �]�N�0�$G�I�}$�1 ���1�0�A L���F�}$F�ERFN� M�NcF]I�J�TANCb �,�J RǱ �^�$JOINT,������3M� �Q���FECE�q��S��bp(D���Q�k �pUS�?��LOCK_FO�`�[�� BGLV��GuLXT  _XM`�AEMP�@�� -P<B2�@$US�!�0"p2*��4QQRW�8�@QQ�SCEj�CNrP $K��M#TPDRA�0�T�A�VEClp�V�@IU�QQVQHE�@TO�OL�s�SV�tREN�PIS3|s�T64�N)`ACH� ���Q3ON��$29�"�P�I�  @$R�AIL_BOXEz���ROBO"T;?�r1HOWc>d<� aROLM�"ge�_�
dxb��/`�p6�O�_F��! � �2�Q^q�N P+�R�PO]r�B�p<�A�`  d�3~	X2MU�֡���@	 IP#VNK��R/b��Q
�QQ�`�PCORDED�@���`b�' |��S1 D )0OB�٣�@dwSq�#pE Sr�ۡSYSSq�ADR =QTCH>��  , �A�A_D�th�*�{Mx�VWVA�� � �P�2kPREV_RT���$EDIT�V/SHWR����$��K��IND� `;�$��D&�[�U�6��KE��� ��l�JMPppLj��TRACE)�[p�I,PSڢC� �NE�Pۡ��TISCK�S��Mo��q���HNR1 @]p��L	_GK&f��gSTY�aLOD1�, �����~� tk 

 G�u%$�q�D=� SFp!$@��8��!�F �P���LSQUaLO<���TERC� ݱ���TSz� @h0�� p��㡼Qb,�O� �#dIZ4$A��! C�"!��oUTPU��1�_�DObB�pXS�@KNjAXIP��cVQcUR���0i#$TH`��~vK���_�P�rEET��P Rlp��O��F��P�A������$ cc>   zÑR3� lѐ u��a��������� ���ù�ӹR���R� �R��d�~�B�d���$�҂�C翐�C���p �2�D�Y�SSC,0� ! h�0DSh�� X}�AT���<�� ~���"ADD�RES�SB�SH�IF�HP_2CH�� zqIK0���T�XSCREEUr"z	 k�TINA�3x@��D �`sQ_��T0# T�� �0'�g00�^��r^�|�RROR_vA���(�h$  ��UE5$$ ��Щq09S�1�qRSM��T�UNEX��j���S_�3��G�ѽ����G�C�B��� �1# 
z��%�="�2��MT!�L�v�m�w0O�D��UI_� HP� O& 8e�w@_T���f� R���Bcg��"�R�O��T0'����7$BUT�T��R RraLUM���u���ERV��R�Pa@��S1({ ^ƠGEUR&SF����A)� LP���E��C�)#�S�1�c�1�T�P0�5.�6.�7.�8����a@����%�Q�AS�'�R�USR�4) I<Z0� UB�AI΀�@FOC�Q@PR�IΡm`�� TR�IP�m�UN$ 5$*	@t�$ k�cj��HR���� �+a��� �G `\��1���\OS��qR��V�H�QS1,`�?�3�>��tH	U�S1-������HOFF!PT0.�[p�O' 1�,�09-�0GUN_WIDTH��>�B_SUB�"p0N�SRT� �/���vA�` �OR`�R�AU��T�����VCC�М�0 ��aC36MFB1�24 ��/0.D1�h %bTq�� �4.��c)�C�`	%�DRIV���_�Vu�,$(��@D��MY_UBY��$V� vA�� B�tC�#�QtB�i0pp+��"L7�BMv�1$��DEY!��EXG�n��Q_MU��X�10orbҲ�}GðPACIN΁}�RGC�52�20�32���!RE{�����Q����2�02^�TARG�@P1R�c0 �R� �03s d��_�FLA΀�r	�"N�RE�#SW0_A1 �@�!�O���A���3��E��UB�a ��HKG�4����:� ��05�!CEA���+GWOR!P�5 �\�MRCV�5� ���OS�M!PC�2S	hB`3hBREFF�FqF\A�0�࿣ �0��mJ�A~J�A�K�EqFO_RC,KXEK�V�S���']#�6�9��6 �$����1؄��b%�pROU��[2�# 1z52�2�P$���� �F΀3��2���Kq�7SUL��4;r��6�5� �P@�3�c�N�f��f��c�PL��#5e�#5e��Ag����$��70 &(��ǡ4� ��C�`+�LO�A�d�a� �iu���`ܓC�pMI��F�R�hTj��fR[$H�Oh��r�`COMM'#��OB�v{X���؇VP]2�HqO_SZ3cQu6/cQu12��Nx0Lx�`�LxWA�eMP�zF�AI�`GT�`AyD�y�!IMRE~T�r_�GP��� ���&ASYNBUF�&VRTD���q6σOL��D_�:�uW�P�ETU�#�`Q�0�ECCUP8VEM:0�e���gOVIRC�q2�Lle��8^Q�0CKLA�S^	�VLEX���9/���l��	�LDLDE��FI<� �r����E���Tp�Q��:����T1�'��β��V�� ;�`��L���{,�"UR�3�0_R�p󔟑�! ���U3�/�/�$�`70���0Ғ �TI�Q��'SCO�� �Cz�4 ;#6;�;�;!� ;/�//%*ᢕ����D�SЧ@ |_�M<)����J*��%��q�=8)G�eLIN�Л�W�@XSGAq�>�  ��N�BPK�cH��HOL�� ���ZABC}?�v2`�XS�@
 |��ZMPCF}@�<�������l!LN�I�΀
��� ~A� ���q+@��CM�CM0CKsCAR�T_ٱ#�P_�� $J����������S��S��2UsXW� ��UXE�!A�<��9��d�J��\�J�l� T�ZPץB ��bOBդ��Y!�D" �Ca⣖�IGH�&3G�?(!�!��A�\���D � �T��A~�$B�PK��'3PK_a�	c�R�V�`F��Ba�OVCY����TU�O0��Jj�
RI��1uD��_TRACEx�V
1}��SPHER��E ,!��������L�$Tb� 2������� d ���? �	 _HD)̀� (���0�fff(�C��nA)�K�Z�$�6��APZ�\�n������q�A�Ȣ���C�p�9�	�=�A��B�������!�3� E���c�����@y�� ���������&C� n��p�  �	V3.0�0�	r85lN�	*� ����B�� ?L��?W�33�x��p	� �  � ?���Cz��_f�x��  ������� �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?O��	  O2OO^OlI0pO�O DlO�O�Kz�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bO>O�JO���O ��O�(��O0�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯t���.��@B��v������J��7 �� Vf���2f������	 2?�*�c�Nχ�rϫ� �ϻ��������)�� M�8�q�\�nߧߒ��� ���������#�I�4�m�X��|������ ��������8�#�\� G���k����������� ����"XC| ���I�s���� �!E3UWi �������� /A///e/S/�/w/�/ �/�/�/�/?�/+?? O?a?k��p?�?�?>? �?�?�?�?�?OOBO 0OfOxO�O�OZO�O�O �O�O�O_,_>_�O
_ t_b_�_�_�_�_�_�_ �_oo:o(o^oLo�o po�o�o�o�o�o �o $H6X~l� ������?�&� �?�h�V���z����� ���ԏ
��.���� d�R���v�����П� �������*�`�N� ��r�����̯��ܯ� �&��J�8�n�\�~� ����ȿ���ڿ��� 4�"�D�j�Xώ��:� ����tϢ�����0�� T�B�x�fߜ߮����� ���������P�b� t��@�������� �����L�:�p�^� ��������������  6$ZHjl~ ������ 2 ��J\n��� ����/
/@/R/ d/v/4/�/�/�/�/�/ �/??�/<?*?L?r? `?�?�?�?�?�?�?�? �?O8O&O\OJO�OnO �O�O�O�O�O�O�O"_ _F_4_V_X_j_�_�_ �_�_p�_ o�_�_Bo 0ofoTo�oxo�o�o�o �o�o�o,<b P����v�� ��(��8�^�L��� p�����ʏ��ڏ܏� $��H�6�l�Z���~� ��Ɵ���؟���2�  �B�h�o������N� ԯ¯����.��R� @�v�������j�п�� ����*�<�N��^� `�rϨϖ��Ϻ����� ��$�J�8�n�\ߒ� �߶ߤ���������� 4�"�X�F�|�j��� �����������$�6� ��V�x�f��������� ������,>��N�Pb����  9� � �����$TBJOP�_GRP 2W���� ?�/��CH�	�E�� �����X��y�^ �,X�o @� ?��ߐD)̴C2?
C랔���333�����<^�%C��n�?fff?�=q�?L��A�  �A��(/����������ff<��7� d?����?��Ü!A� p/�/B/�v/x/���\�"� ?�[��B ��/~O?  Cd6���C�p��.�!�5�? ?�R��2 ;���CA�જ& B�60@R?�?b?t?�?N& �9A�1YQ@�2$>����?iO�?�??�O 2 �B!Rx:�2�� �
=�?�O Y�O
_ Y4__,_Z_ �_f_ _�_�_�_�_�_ o�_�_:oTo>oLozo��o~D���  �0 5	V3.0}01r85l��*�`���B���o  F��� F�� F��� G� G@ G;� GZ.p�z  G�� G�� G�� G�� G�x G��� H� H�L H'� H�7� HG8 H�V�s�� xr�_� F�0/sFp� ( G3� G�mpG^�?s%pG��6p�� G�\ �G�� G�` �G��[sR =u=+�l�!�!�@j����
��A��oK�y� `�\�n����G����ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤߪ y���߬߮  !p���(�:���^�p� �����	����� �j�)�����u�?� ���������������� ��);M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?OO+O=OOOaO sO�O���߳O��S��O __�O�OK_]_o_�_ �_�_��_����_1� Y�#og�y�ko}o�o�o �o�o�o�o�o1 CUgy���� ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i��O�O���O 7_տ�����Ϳ/�A� S�e�wω��_���_�_������$TCPP�ACTSW  ^e����IR e��#�CH  ��SPEED �2� C�e�  ��î��_CF/G 	2�#Ѵ����!Ү��_S�PD��
�>�  ��Q#�:�o®��������NU�Mд���
��OU�T 2��
   ����t��n���� ����������/�"�S��F�X�j�|��ZERO��  ���F�ESTPARS��#����HR��AB_LE 1����R���ٔ�����Q���Ѯ���	���
����������4���RDI��<�&8J\�O����H0��S��� �
 �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?����� z�w���Yk}������n2/� *2�P`�0 3�4�L���2�A@���`�IMEBF_�TT���5��&ќCV�ER2�!ѯF�ќ@R7 1�8�0�:� ��H�7a�6����O�1S�� DP �[°�,_���� �0[}��__��)�� ���^Ĕ_�Y?�+�~P3�^��_k�QR[�oo(o1�<oNo`o�to�o�oɬo���|	���`_�$_����ɟ�oV��o��ʿ��8V�T�ox1͌��������V����SS���T�4��yR�bT�l�x���Ҥ�"��X3�Ə���܏�� ���� 0�B�T�GkUh�z�T�7�8����"��O�؟��T�M�@�#�U�N q?H�Z�T�� 䀯��T������ʯT�0P���T���o9��K� �`�r���L@.���E��A.�!�@��� �MI_CHA�N�G 
�DBGL�VͰ�E���ET�HERAD ?j��i����0r��:eu�4:13:�c7:da r�b(��5���dP�RP��@!��!�����~�SNMASK^����o�255.�$�0��#�5�G߁�O�OLOFS_DI����L�ORQCT�RL �ɦ3�:��5�T������� �0�B�T�f�x��� ���������������;�*�_���PE_D�ETAI<ȉָAP�GL_CONFI�G WIgA�?�/cell/$�CID$/grp1�\�c�����
*����2(]o���4��3��� )���40e w���<���� �/ /2/�V/h/z/ �/�/�/?/�/�/�/
? ?.?�/�/d?v?�?�?�?�?*��}S?�?OpO*O<ONO  O�uOTN�R?�O�O�O�O �O_L?)_;_M___q_ �__�_�_�_�_�_o o�_7oIo[omoo�o  o�o�o�o�o�o�o 3EWi{��. �������A� S�e�w�����*���я �����+���O�a� s�������8�͟ߟ� ��'���K�]�o���𓯥�����U�ser View� ��}}1234?567890��� ��0�B�J�Ӱ��j���ΩK	�?����Ͽ��� e�w�բ�	 ��_�qσϕϧϹ�� *ψ�SN��%�7�I� [�m����ψ�5�ϼ� ��������u�7�}�6��p�������)���}�7_�$�6�H�@Z�l�~����}�8� ������ 2��S�Y lCamera٪���@������BE� .@�Zl~�����  r��� //(/:/L/^/�/ �/�/��/�/�/ ??$?K�rBɻ/p?�? �?�?�?�?q/�? OO ]?6OHOZOlO~O�O7? I7��'O�O�O __$_ 6_�?Z_l_~_�O�_�_ �_�_�_�_�OI7��_ Jo\ono�o�o�oK_�o �o�o7o"4FX jos^��o��� ����o2�D�V�� z�������ԏ{I7 �k� �2�D�V�h�z� !���������
� �.�@��I7��ן�� ����¯ԯ母�
�� .�y�R�d�v�������S�e�98�����#� 5�G��X�}Ϗ�6��π���������߮�	t0��Z�l�~ߐߢ� ��[������ߣ� �2� D�V�h�z�!�3�y { �������	��-��� Q�c�u���������� ������t���?Q cu��@���� ,);M_ @�S;������ /�)/;/M/�q/�/ �/�/�/�/r��Kb/ ?)?;?M?_?q?/�? �?�??�?�?OO%O 7O�/�+k�?�O�O�O �O�O�O�?__%_pO I_[_m__�_�_JO� �{:_�_oo%o7oIo �Omoo�o�_�o�o�o��o�o�]   �Y>Pbt��������   }y?�ƓB�  *��]>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h��z�(x  
�`( � �2p( 	 �������ο�� (��8�:�Lς�pϦ����ϐ�z � ^o�!�3ߦoW�i�{� �ߟ߱߸S�������� F�#�5�G�Y�k�}��� ������������ 1�C���g�y������ ��������	P�b�? Qc������� �()pM_ q������� 6/%/7/I/[/m/� ��/�/�//�/�/? !?3?E?�/i?{?�?�/ �?�?�?�?�?OR?/O AOSO�?wO�O�O�O�O �OO*O__+_rOO_ a_s_�_�_�_�O�_�_ �_8_o'o9oKo]ooo �_�o�o�o�_�o�o�o #5|o�ok}� �o������T 1�C�U��y������� ��ӏ���	��b�?��Q�c�u���������@� ��ȟڟ쟻������)frh�:\tpgl\r�obots\r2�000ib&�_185l.xml�� P�b�t���������ί����� �dummy"�;�?�Q�c� u���������Ͽ�� 
��.�;�M�_�qσ� �ϧϹ��������� *�7�I�[�m�ߑߣ� ������������� )�;�M�_�q���� �����������%�7� I�[�m���������� ������!3EW i{������� �/ASew���������;� �88�?��"/� /@/B/T/v/�/�/�/ �/�/�/?�/?B?,?�N?x?b?�?�?�;�$�TPGL_OUT?PUT ��_  � �?O���3;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_�_�3 �@2345678901�_ �_�_�_o o(c��_ Ooaoso�o�o�oAo�o@�o�o'�j}1 Yk}��9K� ����1��?�g� y�������G������ 	��-�ŏ׏c�u��� ������U�˟��� )�;�ӟI�q������� ��Q�c����%�7� I��W��������ǿ _�տ���!�3�E�ݿ �{ύϟϱ�����m� ����/�A�S���a߀�ߛ߭߿���i�A} !��+�=�O�a�r��@/���* ( 	 �_����� ��%��I�7�Y�[�m� �������������� E3iW�{� �����/�V� "7ewS� �����RP
// �@/R/0/v/�/��/ �/`/�/�/�/�/*?<? �/`?r??�?�?�?�? �?H?�?O�?OJO\O :O�O�O�?�O�OjO�O �O�O"_4_�O _j_|_ _�_�_�_�_�_R_o o�_BoTo2odo�o�_ o�o�oto�o�o, >�obt��� ��J\�(��L� ^�<��������ʏl� ڏ �ޏ��6�H���l� ~� �������؟�T� �� ��V�h�F��� ���¯ԯv���
�� .�@���,�v���*���྿��������$T�POFF_LIM� K|�ӱ��|��N_SV��  x�%� ��P_MON �CG�*�|�2�x��STRTCHOK CE���M�VTCOMPA�T:���I�VWVA/R Z���h�K�� ��|�m���_DEFPR�OG %��%�FOLGE011�ߢ�_DISPL�AY���/�INST_MSK  ��� k�INUSsER��-�LCK�����QUICKMEyN��q�SCRE��C��t_scq���!�&�%�7��ST��E�RACE_CFG Z�����	�
?����HNL 2"��#���� ��� �����"�4�F�X�j����ITEM 2��� �%$12�34567890<����  =<����<����  !�����Jӫ�k�� ���);_ �/U���� 	�7�	// ?/���A/��/�/ �/3/�/W/i/{/�/M? �/q?�?�/�???�? A?Oe?%O7O�?MO�? O�O�?�OO�O�O�O aO	_�O�O�O#_�Oy_ �_�__�_9_K_]_�_ �_�_Soeo�_qo�_�_ �o#o�oGo}o/ �o�o|�o��o�� SCUg���� [���������-�?� ��c��5�G���S�Ϗ ��w�ş)����_� �����^���y�ݟ�� ���ů7����m�-� ��=�c�u�ٯ����� !���E���)ύ�M� ��ÿտY�q������ A���e�w�@ߛ�[߿� ߑ��ϧ��+��߀��S����F�� 3 u�F� ��P�F�
 ]��j��~(�UD1:\������R_GRP� 1 ��� 	 @P������@1��U�C�y�g���� ����s����������?�  )I 7m[���� ���3!WEg�	�ա�q� �m�/�'//7/]/ ���/���/���/� k�/#??G?5?k?Y? �?}?�?�?�?�?�?O �?1OOAO���O� �Oe/�O�O�O	_�O-_ k/Q_�/x_�/u_�_QO �_MO�_�_oo'oMo ;oqo_o�o�o�o�o�o �o�o7uOSe #_�_����� �M_3��_Z��_~��_ ����ՏÏ���� �A�/�Q�S�e����� �����џ�Eo5��G��SCB 2!� �����������ϯ������X�_SCREEN �1"��
 �}�ipnl/X�gen.htm$�w���𛿭���P�Pa�nel setu�pü}	index.STMÿ���1�C�U�̷
Rob�ot Info e�9�ϱ��������� �τ�1�C�U� g�yߋ�߯�&����� ��	��-�߶�c�u� �����4�b�X�� �)�;�M�_������ ����������x��� 7I[m�6 ,���!3��W3�UALRM_�MSG ?D��Q� RD��� ���/
//:/@/�q/d/�/�/�/mSEoV  {�&�kECFG $Ne�  D7�A1�   B�Nh�\Q�0�4�  �A 6aX�\��2?=\X�r�~J?7�X�s'b?�3uX�v8�d>��X�}|�?/�X��?9�X�����?6�X����?+�X�T�~�?.�X�[O�!�GRP 2%e�� 0*21�p>�f�j�_f�?�
���a��I�?_g+�/q��O�gO�O�O�O�O�,I_?DEFPROw+F�� (%$UP�023.$_-U00�11  %MA?KRO050�OD%�/_j_�_�_�_�_��_�_o!ooEo�GI�NUSER  �]�ONoI_MENHIST 1&e�  ( P���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,15?3,1 1 �`�o0'D�'�o�o98�`@P,354�ș�:z.HZued�it�bFOLGEpr3���/�:���j37�a25,6�<�������A��oa�381�`24�o�"��4�?�)ԏZ{�,2�D�������E�O�i�9 lq�`��*�<�˟ݟ�m7���������ϯ�6a�a6o��� �2� D�V��s므������� ȿڿi����"�4�F� X��|ώϠϲ����� e�w���0�B�T�f� �ϊߜ߮�������s� ��,�>�P�b���� ����������ݯ� (�:�L�^�p������ �������� ��$6 HZl~��� ����2DV hz����� �
/�./@/R/d/v/ �/�/)/�/�/�/�/? ?�<?N?`?r?�?�? �?�/�?�?�?OO&O �?JO\OnO�O�O�O3O �O�O�O�O_"_4_�O X_j_|_�_�_�_A_�_ �_�_oo0o�_Tofo xo�o�o�o�oOo�o�o ,>)?�ot� �����o��� (�:�L��p������� ��ʏY�k� ��$�6� H�Z��~�������Ɵ ؟g���� �2�D�V� ���������¯ԯ� u�
��.�@�R�d�Oz��$UI_PAN�EDATA 1(�������  	�}�/frh/cgt�p/doubde�v1.stm o�de=1 lse� ave&ACT�ION=101&C2=7p������  )prim�<�  }?�c�u�0�ϙϫϽ� )���� �����+�=�$�a�H� �ߗ�~߻ߢ���������Lv�� �5� 5(nM¦�2��]�o���<���dual���� O� ��$�6�H�Z�� ~�e������������� ��2V=z�s�#������� ,>P�t�� ������Y/ (//L/3/p/�/i/�/ �/�/�/�/ ?�/$??H?Z?-� �_?�?�? �?�?�?�?D?O�9O KO]OoO�O�O�?�O�O �O�O�O_�O#_G_._ k_R_�_�_�_�_�_�_ �_n?�?1oCoUogoyo �o�_�o"O�o�o�o	 -�o?cJ�n �������� ;�"�_�q�X���oo ˏݏ���%�x�I� [��o�������ǟٟ @����!�3��W�>� {���t�����կ��� ��/�����?�w��� ������ѿ$���h�� +�=�O�a�s�ڿ�ϩ� ���ϴ������'�� K�2�o߁�hߥߌ��� ��N�`��#�5�G�Y� k�ߏ�ϳ������� ���t��C�*�g�N� ���������������� ?Q8u��������� )�7��&cu� ���$��/� �;/"/_/F/�/�/|/ �/�/�/�/�/?��������$UI_PO�STYPE  ���� 	� ?v?E2QUI�CKMEN  �T;c?y?G0RESTORE 1)���  �?���?�3�?��mODOVOhOzO�O /O�O�O�O�O�O�O_ ._@_R_d_Oq_�_�_ _�_�_�_oo�_<o No`oro�o�o9o�o�o �o�o�_!3�o n����Y�� ��"��F�X�j�|� ��9C�����1��� �0�B�T���x����� ����c������,� ׏9�K�]�ϟ������ ί௃���(�:�L� ^����������ʿ�7oSCRE�0?�=u1sc�0Wu2�3�4�U5�6�7�8�E2USER����Sks�f�3f�4f�U5f�6f�7f�8f��E0NDO_CFG� *T;� �E0P�DATE P���KS_24��1G�_INFO �1+�����10% пߣ��D�'�h�z� ]ߞ߰ߓ��߷���
���.�@�#�d�}<��O�FFSET .�=q�l��0s����� ������!�N�E�W� ��[��������������/y��?{
�j�}�UFRAM/E  d������RTOL_ABRqT����ENB�~�GRP 1/�9��1Cz  A� :8l�8J\n�B����
�0U����MSK  h���	N�%���%KH/�2VCCMf��0��]"MR {26T9 d�Կ¼�	��O�~?XC56 *�/�&�X�����5���A@�p��L. �8?d�7?@I?v?�!q?�?5�A�l��?�?l�� B����1l��5�? Ob??OOcONO�OrO �O�O�O�O8O�O__ _M_ Oq_�_d��!�! �/�_�/�/�/??'? o�O\oSo1_�o�o�? �?�o�?__�o"io{o =jU�y��� -���	�B�U_f� x�����!�_���_�_ �_oo'o��\�S� 1������o�oڟ�o_� ��"�i�{�=�j�U��� y�����֯-���ɯ� 	�B�U�f�x����=� ����͏ߏ���'� ��\�S�1��ϤϷ� ɟ���_���"�i�{� =�j�Uߎ�y߲ߝ��� -������	�B�U�f��x�O/ISIONT�MOU� $r%����d#7�0 ��1t/ �FR:\��\DA�TA\�� ��� MC��LOG���   UD1���EX��' B@ ��O� �7/m� �q����� �  =	 �1- n6 � -��T�L�&,x�����=������T���TRA�IN6������"8�+ (:���S.� Sas����� ��'9KX&/LEXE��9�+�!�1-eR,MPHA�SE  k%�#��R]!SHIFTM�ENU 1:�+
� <\�6//�����!/Z/1/C/�/g/ y/�/�/�/�/?�/�/�D??-?z?Q?	L�IVE/SNAP�n3vsfliv��?^3�� SE�TU�0�2menu �?�?d?)O;OB��3;����	(H'OЌO\����� ��@Z�A�B8`�`�!������A�B��C簝�G ��KSFMaE�0����� �kMO�<��z���WAITDINE�ND���Q@WOK�  �X[]��w_S܋_^YTIM�����\GH_�]j_�[�_��Z�_�Z�_\XREL�E�gU@T���=�AS_ACT�0
h��a����d�� =���b%$FOLG�E011.	r0�004��dRDI�S�0�oAPV_AX�SRG`2>bJ<��O��Gp4 _IR  ��᥀���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z���ޖ�ZABC31?LbI�� ,�=�2�� ܬ¯�����
��Y����MPCF_G 1@S}0A��������ҿ������,�b�M�P��AbI  ��@���:��Q8�|O����t��Ϙ�?�T�������D���� k�-ߞ߰��ѿp��� ��������	�l�E�� i�{�ߟ�R�\�n߀� �������2���e�w� ���������.� �d�=OZ�s�@� �\�����' 9����Tf���� �&�/5/� \//�/B/T/f/x/ �/�/F��(?:?L?�v>��u�(PBS{j�P�_CYLINDE�R 2CS{ ���& ,(  * �?�=�#�?O�?8OM �/nO�O�N�?�O $O�O�O�O_RO3_E_ W_�O{__�O�_�_�_��_*_oof�R�2DSw�`�P�"�hoxl�s �/�o�o�o��o�o�1�qA��o*yo�o `�o��o}�	� �?y&�uJ��Z� ���m����?��׏��_�4�F����2SPHERE 2E�=�o_���_��͟��� �_L�'�9�i_]���� ��z���������F� X�5���Y�@�R���֯�ſ׿N�ZZ  �$��4