A��*SYSTEM*   V8.2306       4/24/2014 A 
  *SYSTEM*  �MN_MCR_TABLE   � $MACRO_NAME %$PROG_NAME %$EPT_INDEX  $OPEN_ID  $ASSIGN_TYPE  $ASSIGN_ID  $MON_NO  $PREV_SUBTYP  $USER_WORK  $SYS_LEV_MSK  $MCR_RTN  �MN_MCR_SOP_T  � $SOP_EMGOP  $SOP_RESET  $SOP_REMOTE  $SOP_HOLD  $SOP_USER1  $SOP_USER2  $SOP_START  $SOP_PDI8  $SOP_PDI9  $SOP_PDIA  $SOP_PDIB  $SOP_PDIC  $SOP_TPDSC  $SOP_TPREL  �MN_MCR_UOP_T  � $UOP_ESTOP  $UOP_HOLD  $UOP_SFSPD  $UOP_CSTOP  $UOP_RESET  $UOP_START  $UOP_HOME  $UOP_ENBL  $UOP_RSR1  $UOP_RSR2  $UOP_RSR3  $UOP_RSR4  $UOP_RSR5  $UOP_RSR6  $UOP_RSR7  $UOP_RSR8  $UOP_PNSTRB  $UOP_PDSTRT  �$$CLASS  ������       �$MACROLDUIMT         �    �$MACROMAXDRI         �   
�$MACROTABLE 1 ������ � d%Open hand 1                           %ZG_MENUE                              _        s<h   %Close hand 1                          %                                       ��               %CUST_MN nd 1                          %CUST_MN                               �        s3�  %CUST_MN d 2                           %CUST_MN                               �        s1$  %Close hand 2                          %                                       ��               %Relax hand 2                          %                                       ��               %                                      %                                       ��               %                                      %                                       ��               %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %
Send Event                            %SENDEVNT                              =               %	Send Data                             %SENDDATA                              <               %Send SysVar                           %SENDSYSV                              >               %Get Data                              %GETDATA                               ?               %Request Menu                          %REQMENU                               @               %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                %                                      %                                      ��                �$MACRO_MAXNU         ��   ��$MACRSOPENBL �������                                                      �$MACRSPDIMSK      ����    �$MACRSPSUMSK      ����    �$MACRTPDSBEX         �    �$MACRUOPENBL �������                                                                       