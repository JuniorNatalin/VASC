A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DCSS_IOC_T   P $OPERATION  $L_TYP  $L_IDX  $R1_TYP  $R1_IDX  $R2_TYP  $R2_IDX  0�$$CLASS  ������   P    P�$DCSS_IOC 2 ������P @             
                      
                       
                     
                      
                                                   
                  ����                                              ����                                                                            	                  	   
                     
   
                                            ����                     ����                      ����                      ����                    ����   ����   	          ����                        
   	                  
   	                      
                    
                     
   
                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$DCS_C_CCL ?������P  	All param             
Base param            Pos./Speed check      Safe I/O connect      �$DCS_C_CCR ?������P  	All param             
Base param            Pos./Speed check      Safe I/O connect      �$DCS_C_CSI ?������P @ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_CSO ?������P @ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_NSI ?������P   �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_SIR ?������P @ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_SPI ?������P @ SFDI1                 SFDI2                 SFDI3                 SFDI4                 SFDI5                 SFDI6                 SFDI7                 SFDI8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �$DCS_C_SPO ?������P @ SFDO1                 SFDO2                 SFDO3                 SFDO4                 SFDO5                 SFDO6                 SFDO7                 SFDO8                 �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_SSI ?������P  SVOFF                 FENCE                 EXEMG                 �                      NTED                  OPEMG                 AUTO                  T1                    T2                    MCC                   CSBP                  �$DCS_C_SSO ?������P  C_SVOFF               C_FENCE               C_EXEMG               C_SVDISC              C_NTED                C_T1                  C_T2                  