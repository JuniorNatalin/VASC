A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �CELL_GRP_T   � $CELL_FRAME $MOUNT_LOC $CF_METHOD  $CPY_SRC_IDX  $PLATFRM_OFS $PLATFRM_DIM  $BASE_OFFSET $BASE_DIM  $AUX_ORDER   $AUX_XYZ_MAP   $AUX_OFFSET   $AUX_LENGTH   $ATTCH_GP_MS  $AUTORAIL  �$$CLASS  ������   D    D�$CELL_FLOOR         D8�?�              ?�              ?�                  �$CELL_GRP 1 ������D H8  ?�      �       ?�              ?�          D'�     8  ?�      �       ?�              ?�          D'�        ���8�������������������������������������������������8�������������������������������������������������  ���������  ���������  ���������  ���������������8  ?�      �       ?�              ?�                  8!  ?�      �       ?�              ?�                     ���8�������������������������������������������������8�������������������������������������������������  ���������  ���������  ���������  ���������������8  ?�      �       ?�              ?�                  81  ?�      �       ?�              ?�                     ���8�������������������������������������������������8�������������������������������������������������  ���������  ���������  ���������  ���������������8  ?�      �       ?�              ?�                  8A  ?�      �       ?�              ?�                     ���8�������������������������������������������������8�������������������������������������������������  ���������  ���������  ���������  ����������������$MNUFRAME A������D d  88�?g�,�ڐ/;{��>ڍ?g�?;��K��Wݻi�&?�nE,��D����>�    8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                    88!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                    881�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                    88A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  �$MNUFRAMENUM      >   D      �$MNUTOOL A������D \  88�?�          �   ?�          �   ?�          D�Ff    8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                    88!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  8!�?�              ?�              ?�                    881�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                  81�?�              ?�              ?�                    88A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  �$MNUTOOLNUM        D  