��   ɋ�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_CPC_�T   � �$COMMENT� $ENA�BLE  $�MODJGRP_�NUMKL\ � $UFRM�\] _VTX �M �   $Y��Z1K $Z2��STOP_TY}PKDSBIO��IDXKENBL?_CALMD�&}S. � 8�J\TC�u
SPD_LI_����COL�&Y0 � � !CHG�_SIZ$A�P7ECDIS � � �7�C�����Jp 	�J �� ��"��$�'"_SEs�DxSTAT/� D $FP_�BASE �$LINK`$!��j&_Vs.Hs# ��&J- ���ZAXS\UPR:LW�'CU�� Ԡ$� | 
�/�/�/4�??j�&ELE�M/ T $1Uc c1j"NO�7�0�a3UTOOi�2H�A�4�� $DA;TA" �4e�0   @P:�0 _2 
&PP%' ��P!U*n   oFSyCjrB�� zB(�F�D(�1R|5C�DROBOT�H��CQBo�E�F$�CUR_"�BH$SwETU�	 l� ��P_MGN�I?NP_ASS�  @�� �3�8"7GP U��>VhSP!��&T1�
@B\8�8�T= �0 P�+ Kec1V�RFY�8�T$5&1ȕ ��W��1$�R�|TPH/ ([ �#A�#A��#A3tBOX/ 8�0������`bo%c�TUIR>�0  ,[ �6�2`ERa02 �$k` �a_mS�bX�fZN/ 0 [9&0� �arZ_� �_p� tu0  @�A��Yv	�on��$�$CL,P  �����q��Q��Q��$' 2 �u�Q   �Q�q���b0�p
�}�p��~�4� F���m������ ǏُL�������E� ��i�{���$�6� �Z�����A���Ɵ ؟��������2��V� h�z�+���O�a�ԯ�� ��
�@�Ϳ����v� 'Ϛ����п^ϓϥ� ���<�N���r��5� Gߺ�k����ϡ���� ����\��ߒ�C�� g�y��ߊ��"�4��� X�	����?������� �������0���T�f� x�)��M_����� �>�t% ���m\�� �:L�p�3/E/ �i/��q//�/�/ �/Z/?~/�/A?�/e? w?�?�/�? ?2?�?V? OO�?*OOO�?�?�O �?�O�O.O�OROdOvO '_�OK_]_�O�_�O_ _�_<_�_�_r_#o�_ �_�_ko�_�o�oo�o 8oJo�o�o1C�o g�o�o"��� X	�|���O�u� ������0��T�� �)���M���ҏ���� ����,�ʟ�b�t�%� ��I�[�Ο���� ǯ:����p�!��������i�ܯ������$�DCSS_CSC� 2I�ɱQ  D�� �@���&���J�\� n�=ϒϤ϶υ����� ����"�4��X�j�|� Kߠ߲��ߓ������ ��0�B��f�x��Y� ������������� >�P�b�1�����g������������GRPw 2ɻ ��	��cN�r� �����; &Kq\���� ��/�%//I/4/ m/X/j/�/�/�/�/�/ �/?�/3??W?B?{? f?�?�?�?�?�?�?�? OOAO,OeOPO�O�O �O|O�O�O�O�O__ _O_:_s_�_T_f_�_ �_�_�_o�_'oo7o ]ooo>o�o~o�o�o�o��o�o�o5
S?TAT 2ɹY��,8���k>�6?L��?
X_�+���?�!?���?:��>��;rC��:Ce?�PEn�ɱ,p�8xq?h�>��^\��q+4���?�  �q���p4��ZC��b�C��p  �ɱxr1�5����`?$�@�$������D�6�y�����X�%�D,�b�vH�����`c? �)��^a�p��=Ѿ�b��Xb'�]���� 
&Õ>��DH���u����Q�">ѷՈ@�jD�H��?�K��Q�����[B�v(Bj��E�G�u�=~���;9�?f��K��?Q�>��X���¿:����;x��z�� ́ɵ��ɵ�J�\� :������z�r���� �uğ�؟�$�� � B�D�V�x�������د �w���d��H�Z�8� ~�����䯺���ƿ� ڿ��&��2�\�F�h� ��|ώ��ϲ�p�
�߀��@�R�0�v߈�f�>��lk�d�޽��s�ZƟ��˯뾪�V>���K>W�ѿ�p�XDK�C�}D����zvG�>��U)q����[4�"X��r�п���r���B�N��zUH���r�?  ����H����]�������=�(�jD`��X�࿱���M?c�����^��ߴ�n���[&�x�����F�-�L�D�D8n,X��̑��O?Wa�ol�p�t��E>�替p�����D<�CU{"D�����gԷ>����>�~O�����?p�=������B�W��?p�Z��߸� ��l�>�P�.�t���d� �������������� (R<N�r� ������6H ��l~\���� ��/�/2/4/ F/h/�/|/�/�/�/�/ �/$.?@?�d?v?T? �?�?�?��������� ��&�8�J�\�n�� �����������?�? "��?n_�?^_�_�_�_ �_�_�?o�/"oLo 6oXo�olo�o�o�o�o �o�o�o$�_fx V������_8 ��D�.�P�z�d� v�������ΏЏ�� .��^�p�������� ʟܟ�?,_>_�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__�� R_��������Կ��� 
���<�F��R�|� fψϲϜϾ������� ��*�T�>�ϖ�� �����߼���.�h� >�D�J�t�^���� ��������� ��L� 6��ߎ���~������� ����\�n�,�>�P� b�t���������ί� ���(�:�$6H �������/�(/ :/ �J�d/n�`/�/�/ �/�/�/�/�/??$? N?8?Z?�?v��?�?/ �?�?�?O2OL/^/�? nOt?zO�O�O�O�O�O �O_�O_F_0_R_|_ f_DO�_O�_�_o�_ *o<oz��\n� ������� "lFXjTofoxo o���"�4��X� j�PO�_���_��ʏ�� Ə ����� �2�T� ~�h������_���H� �,�
�P�b�|����� ʟ���������
��� �@�*�L�v�`����� ҟܿ�@���$��4� Z�8Ϫ���o�o�o �o�o�o�o
.@ Rdv��߄ϖ�� J��.��R�d�B�� ���������� �0��<�f�P�b��� ��������z�& J\:������� ������($ FHZ|���� //pB/T/2/x/ �/t����ߪϼ����� ����(�:�L�^�p� �ߔߦ߸��ߴ/�/ � �/LO�/\O�O`OrO�O �O���O� _*__ 6_`_J_l_�_�_�_�_ �_�_o�_�ODoVo4o zo�ojo�o�o�Oo�o �_�o".XBd �x������ �o<�N�,�r���b�������e�$DCSS?_JPC 2�2�a�Q ( D��%��$�6� H��l�~���_���Ɵ �������ݟ2�D�V� %�z�����m�¯ԯ� ��
�����R�d�3� ������{�п���ÿ �*����`�r�Aϖ� �Ϻω��������&� 8�J��n߀�O�a߶� �ߗ��������4�F� X�'�|��]�o����� ��������B�T�f� 5�������}������� ��,��PbtC �������� (:	^p�Q� ���� //�6/ H//)/~/�/_/�/�/ �/�/�/? ?�/D?V?P%?7?#�؅S���@BS HA�LT�?u5u?  >)�=��ʹ?�?B�4�?�?O�6 O2ODO�6`OrO�O�6 �A�O�O�O�3�O�O�C_�6 _2_�_�6�`_r_�_�6	�_�P� �_ox?$��_Eoo*o {oNo�oro�o�o�o�o �o�o�oA&wJ \n������ �=��a�4���X�j� ����ɏ���֏�9� ��0���T�f����� ������ҟ�"�G�� ,�}�P���t�ů���� ��ί	��C��(�y� L�^�p���������ʿ ܿ�?��$�bχ�Z� lϽϐ��ϴ�����π;��I�2߃�Vߊ?_�MODEL 2Σ;xt�i�
 U<m�c�:�H�J "����X�/�A�S�e� w����������� ��+�=���a�s��� ������������g�P ��+�o��� �����L#5 �Yk}��� / ��6///1/C/U/ g/=�/a�/�/?�/ �/D??-???�?c?u? �?�?�?�?�?�?�?@O O)OvOMO_O�O�O�O �O�O�O�O�/�/�/_ _�_�Om__�_�_�_ o�_�_8oo!o3oEo Woio�o�o�o�o�o�o �o�ojAS� ;_M_{��u�� ��+�x�O�a����� ������͏ߏ,��� b�9�K�]�o������� ��ɟ�����p� �Y�k��������ů ׯ$�����l�C�U� ��y���ؿ����ӿ � ��	�V�-�?ό�'�9� K�yϋ�a�����.�� �d�;�M�_�q߃ߕ� �߹��������%� 7�I��m������ ���&��������E� W���{����������� ����X/A�e w������ B+=��7�e w���/�/P/ '/9/K/�/o/�/�/�/ �/?�/�/�/L?#?5? �?Y?k?�?�?�?�?� O��?�?ZO1OCO�O gOyO�O�O�O�O_�O �OD__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o�?�o#OQoco�o �o�o�o�o% 7�[m���� ���8��!�n�E� W�i�{�����uo���o ǏُF��/�|�S�e� w�ğ������џ�0� ��+�x�O�a����� ��䯻�ͯ߯,��� ����=�O���7��� ��ɿۿ�:��#�p� G�Y�k�}Ϗϡ����� ��$�����1�C�U� ��yߋ���s������� 2���-�?�Q�c�� ������������� �d�;�M���q����� ��������N�� ��);�#��� ��&�\3E W�{����/ ��/X///A/�/e/ w/�/_q��/�/�/ ??f?=?O?�?s?�? �?�?�?�?O�?OPO 'O9OKO]OoO�O�O�O��O_�O�O�O�$�$�DCSS_PST�AT ����cQQ  �  t_�Z r_ (�_�_�WkPkP��_�_ l cdP��P;_4oFo�)�"ocUcUdovoTTSETUP 	cY'B�&T�#�!�d�OYT1SC 2
4�j`�!Cz�#�/}�eCP R�l�� DSoz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ��.h%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� ����������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G����� }��������������� 1CUgy� ������	 -?Qcu��� ����Z�D�/*/ </�/`/r/�/S/�/�/ �/�/�/??�/8?J? ?[?�?�?a?�?�?�? �?�?O"O�?FOXOjO 9O�O�O/}O�O�OoO __0_�OT_f_x_G_ �_�_�_�_�_�_�_o ,o>ooboto�oUo�o �o�o�o�o�o: L�O)���� �� ��$��H�Z� l�;�����q���؏� ��� �2��V�h�z� I����������_ ՟.�@�ǟd�v���W� ����Я������� <�N��_�����e��� ̿޿����&���J��\�n�=ϒϤ�s��$�DCSS_TCP�MAP  ������Q� @ ~�~�R~�~���~�~��~�~�	g�  U~�~�~�~�U~�~�~�~�U~�~�~�~��~�~�~�~��~�~�~�~��~� ~�!~�"~�#�~�$~�%~�&~�'�~�(~�)~�*~�+�~�,~�-~�.~�/�~�0~�1~�2~�3�~�4~�5~�6~�7�~�8~�9~�:~�;�~�<~�=~�>~�?�~�@��UIRO �2����� $��"�4�F�X�j�|� ������������� �0�B�T�}��}� ������������ 1CUgy�� ���^�����- ?Qcu���� ���//)/;/M/ _/��/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?v/�O��UIZN 2]��	 ����� PObOtOy�KO�O�O�O �O�O�O_�O0_B_T_ _x_�_�_k_�_�_�_ �_�_o,o�_Poboto �oIo�o�o�o�o�o �o:L^-�� �i�����$� 6��Z�l�~�M����� Ə؏�����ݏ2�D��V�O��UFRM R�����џ� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߒ� �߱����������� /�A�S�e�w���� ����������+�=� O�a�s��ߗ������� ����'9K] o������� �#5GYk���x����� �//�B/T///x/ �/e/�/�/�/�/�/�/ ?,??P?b?y��? �?I?�?�?�?OO�? :OLO'OpO�O]O�O�O �O�O�O�O�O$_6__ Z_l_�?�_�_A_�_�_ �_�_o�_2oDooho zoUo�o�o�o�o�o�o �o.	Rd{_� �9������ �<�N�)�r���_��� ����ޏ��ˏ�&�� J�\�sw