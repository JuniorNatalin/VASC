A��*SYSTEM*   V8.2306       4/24/2014 A 	  *SYSTEM*  �CELLSET_T   w$GI_STYSEL_P $GI_STYSEL_T  $GI_STYSEL_I  $GO_STYSEL_P $GO_STYSEL_T  $GO_STYSEL_I  $DO_STYSTR_P $DO_STYSTR_T  $DO_STYSTR_I  $DI_INISTY_P $DI_INISTY_T  $DI_INISTY_I  $UI_START_I  $RSRPNS1_T  $RSRPNS2_T  $RSRPNS3_T  $RSRPNS4_T  $RSRPNS5_T  $RSRPNS6_T  $RSRPNS7_T  $RSRPNS8_T  $PNSTROB_T  $ACKSNO1_T  $ACKSNO2_T  $ACKSNO3_T  $ACKSNO4_T  $ACKSNO5_T  $ACKSNO6_T  $ACKSNO7_T  $ACKSNO8_T  $ACKSTROB_T  $RSRPNS1_I  $RSRPNS2_I  $RSRPNS3_I  $RSRPNS4_I  $RSRPNS5_I  $RSRPNS6_I  $RSRPNS7_I  $RSRPNS8_I  $PNSTROB_I  $PNSGIN_I  $PNSDIN_I  $ACKSNO1_I  $ACKSNO2_I  $ACKSNO3_I  $ACKSNO4_I  $ACKSNO5_I  $ACKSNO6_I  $ACKSNO7_I  $ACKSNO8_I  $SNACK_I  $PNSGOUT_I  $PNSDOUT_I  $DI_OPTNA_P $DI_OPTNA_T  $DI_OPTNA_I  $DI_OPTNB_P $DI_OPTNB_T  $DI_OPTNB_I  $DI_OPTNC_P $DI_OPTNC_T  $DI_OPTNC_I  $GI_DECSN_P $GI_DECSN_T  $GI_DECSN_I  $DI_TRYOUT_P $DI_TRYOUT_T  $DI_TRYOUT_I  $DI_PTHCNT_P $DI_PTHCNT_T  $DI_PTHCNT_I  $DO_INCYCL_P $DO_INCYCL_T  $DO_INCYCL_I  $DO_TASKOK_P $DO_TASKOK_T  $DO_TASKOK_I  $DO_OPTNA_P $DO_OPTNA_T  $DO_OPTNA_I  $DO_OPTNB_P $DO_OPTNB_T  $DO_OPTNB_I  $DO_OPTNC_P $DO_OPTNC_T  $DO_OPTNC_I  $GO_DECSN_P $GO_DECSN_T  $GO_DECSN_I  $DO_INTLCK_P $DO_INTLCK_T  $DO_INTLCK_I  $DO_ISOLAT_P $DO_ISOLAT_T  $DO_ISOLAT_I  $DO_MANSTY_P $DO_MANSTY_T  $DO_MANSTY_I  $GO_PTHSEG_P $GO_PTHSEG_T  $GO_PTHSEG_I  $DO_PTHREQ_P $DO_PTHREQ_T  $DO_PTHREQ_I  $DO_TRYOUT_P $DO_TRYOUT_T  $DO_TRYOUT_I  $DO_HFAULT_P $DO_HFAULT_T  $DO_HFAULT_I  $DO_HALERT_P $DO_HALERT_T  $DO_HALERT_I  $DO_HEARTB_T  $DO_HEARTB_I  $DO_HNDBRK_T  $DO_HNDBRK_I  $DO_PRGABT_T  $DO_PRGABT_I   !d�CLMLIO_T   $TYPE  $INDEX  �$$CLASS  ������       �$CELL_OPTION         �   �$CELL_SETUP  ������Style-Auswahl	           Style Anf./Echo          Style Ack                Style starten                                                                       	   
                                                                Option Bit A             Option Bit B             Option Bit C             Auswahlcode              Tryoutmodus              Bahnseg. weiter          In Zyklus                Aufg OK                  Manuel Opt.Anf.A         Manuel Opt.Anf.B         Manuel Opt.Anf.C         Man. Auswahl Anf         Roboterverrieg.          Robot in Isolate         Man. Zyklusstart         Bahnsegment              Bahnseg.Anf weit         Tryout-Status            	MH Fault:                	MH Alert:                   #  �              �$CLMLIO 1������                                                          �$STYLE_COMNT ?�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �$STYLE_COUNT         ��    �$STYLE_ENAB  �������                                                                                                   �$STYLE_MENU         �   �$STYLE_NAME ?%�������   (%$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              %$********                              