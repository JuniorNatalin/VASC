��   ɋ�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_CPC_�T   � �$COMMENT� $ENA�BLE  $�MODJGRP_�NUMKL\ � $UFRM�\] _VTX �M �   $Y��Z1K $Z2��STOP_TY}PKDSBIO��IDXKENBL?_CALMD�&}S. � 8�J\TC�u
SPD_LI_����COL�&Y0 � � !CHG�_SIZ$A�P7ECDIS � � �7�C�����Jp 	�J �� ��"��$�'"_SEs�,xSTAT/� D $FP_�BASE �$LINK`$!��j&_Vs.Hs# � &J- ���ZAXS\UPR:LW�'CU�� ��$� | 
�/�/�/4??�j<4ELEM/? T $Uc c1�j"NO�7�0a3UT3OOi�2HA�4�~� $DATA"� �&e0 �  @P:�0 2� 
&PP% ɘ�P!U*n   oFSyCjrB� zB)(�F�D(�1R5C�D_ROBOT�H�C�QBo�E�F$CU�R_"�B &SE;TU�	 l� ��P_MGN�INP_ASS� @ �� �3�8"7GP U��>VhSP!��&T1�
@B\8�8�T= 0 �P�+ Kec1VRCFY�8�T$5&1� ��W��1$R�UPH/ (�[ �#A�#A�#A3�tBOX/ 8 �0�����`bo�%jTUIR�0 � ,[ �62`ER�a02 $k` ��a_S�b�L�fZN/ 0# [9&0� arZ_� �_� tu0  @�A�Yv	�o�n��$$CL�,P  ���t�q��Q��Q�$'� 2 �uQ?   ��q�J��b0�p�}P��~�4�F��� m������ǏُL� ������E���i�{� ��$�6��Z�� ���A���Ɵ؟���� ����2��V�h�z�+� ��O�a�ԯ����
�@� Ϳ����v�'Ϛ��� �п^ϓϥ����<� N���r��5�Gߺ�k� ���ϡ��������\� �ߒ�C��g�y��� ���"�4���X�	�� ��?����������� ��0���T�f�x�)�� M_������ >�t%��� m\���:L �p�3/E/�i/� �q//�/�/�/Z/? ~/�/A?�/e?w?�?�/ �? ?2?�?V?OO�? *OOO�?�?�O�?�O�O .O�OROdOvO'_�OK_ ]_�O�_�O__�_<_ �_�_r_#o�_�_�_ko �_�o�oo�o8oJo�o �o1C�og�o�o "���X	�| ���O�u������ �0��T���)��� M���ҏ��������,� ʟ�b�t�%���I�[� Ο����ǯ:�� ��p�!�������i�ܯ�������$DCS�S_CSC 2�I�ɱQ  D���@�� �&���J�\�n�=ϒ� �϶υ���������"� 4��X�j�|�Kߠ߲� �ߓ��������0�B� �f�x��Y������ ��������>�P�b� 1�����g������������GRP 2Nɻ ��	�� cN�r���� ��;&Kq \������/ �%//I/4/m/X/j/ �/�/�/�/�/�/?�/ 3??W?B?{?f?�?�? �?�?�?�?�?OOAO ,OeOPO�O�O�O|O�O �O�O�O___O_:_ s_�_T_f_�_�_�_�_ o�_'oo7o]ooo>o �o~o�o�o�o�o�o��o5
STAT� 2ɹY�,8���T�ܽ���6��F���� ?~�]��k��?����~2�U�D�t�-?jD�L�ɱ,p8xq?��:2�N���k{�4��W/?�  �q��p�p�ZC���>Y����ɱxr0-����$?9�߿9�ܺ���p���y������P�DB���u����Q��P?��2�_�q��������2�6(�����º���[D{�;��u;�ٔ��;@�@�3�GH��1�D�p����%DT�A�?�VD}����vU��f�/���:1ԯ��p�:뾠�8��8?�q��{ ��~́ɵ��ɵ� J�\�:������z�p� ����uğ�؟�$� � �B�D�V�x����� ��د�w���d��H� Z�8�~�����䯺��� ƿ�ڿ��&��2�\� F�hϒ�|ώ��ϲ�p� 
����@�R�0�v߈�|f�Ѐr���؀�2���X?~����k�����ו�}���p>?�K��p�|�:wC�3�r��6�v����p��t�>nK}��|����p}��p���p�������۾��?�DB� ���䶳��0�C��{��<��@��C��T�KL������pT��X��w�g��h�o�t��B�s�p���:$��V?"���������uY����:B�޾�p�:K����/8�������� ����l�>�P�.�t��� d��������������� (R<N�r �������6 H��l~\���� ��/�/2/ 4/F/h/�/|/�/�/�/ �/�/$.?@?�d?v? T?�?�?�?������� ����&�8�J�\�n� ������������? �?"��?n_�?^_�_�_ �_�_�_�?o�/"o Lo6oXo�olo�o�o�o �o�o�o�o$�_f xV������_ 8��D�.�P�z� d�v�������ΏЏ� �.��^�p������ ��ʟܟ�?,_>_�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__� �R_��������Կ�� �
���<�F��R� |�fψϲϜϾ����� ����*�T�>�ϖ� 迆����߼���.� h�>�D�J�t�^��� ���������� �� L�6��ߎ���~����� ������\�n�,�>� P�b�t���������ί ����(�:�$6 H�������/� (/:/ �J�d/n�`/�/ �/�/�/�/�/�/?? $?N?8?Z?�?v��?�? /�?�?�?O2OL/^/ �?nOt?zO�O�O�O�O �O�O_�O_F_0_R_ |_f_DO�_O�_�_o �_*o<oz��\n �������� "lFXjTofo xoo���"�4�� X�j�PO�_���_��ʏ ��Ə ����� �2� T�~�h������_��� H��,�
�P�b�|��� ��ʟ���������
� ���@�*�L�v�`��� ��ҟܿ�@���$�� 4�Z�8Ϫ���o�o �o�o�o�o�o
. @Rdv��߄ϖ� �J��.��R�d�B� ��������� ���0��<�f�P�b� ����������z�& J\:������ �������( $FHZ|��� �//pB/T/2/ x/�/t����ߪϼ��� ������(�:�L�^� p߂ߔߦ߸��ߴ/�/  �/LO�/\O�O`OrO �O�O���O� _*_ _6_`_J_l_�_�_�_ �_�_�_o�_�ODoVo 4ozo�ojo�o�o�Oo �o�_�o".XB d�x����� ��o<�N�,�r���b�������e�$DCS�S_JPC 2��eQ (# D��%��$� 6�H��l�~���_��� Ɵ�������ݟ2�D� V�%�z�����m�¯ԯ 毵�
�����R�d� 3�������{�п��� ÿ�*����`�r�A� �ϨϺω�������� &�8�J��n߀�O�a� ���ߗ��������4� F�X�'�|��]�o��� ���������B�T� f�5�������}����� ����,��Pbt C������� �(:	^p�Q ����� //� 6/H//)/~/�/_/�/ �/�/�/�/? ?�/D?�V?%?7?#�؅S���@BS H�ALT�?u5u?  })�=��ʹ?��?�4�?�?O�6 O2ODO�6`OrO�O@�6�A�O�O�O�3�O�OC_�6 _2_�_�6!`_r_�_�6	�_�P��_ox?$��_Eoo *o{oNo�oro�o�o�o �o�o�o�oA&w J\n����� ��=��a�4���X� j�����ɏ���֏� 9���0���T�f��� ��������ҟ�"�G� �,�}�P���t�ů�� ����ί	��C��(� y�L�^�p��������� ʿܿ�?��$�bχ� Z�lϽϐ��ϴ���� ��;��I�2߃�Vߊ?�_MODEL 2��;xt�i�
� <m�c�:�H �J"����X�/�A�S� e�w��������� ����+�=���a�s� ��������������g� P��+�o�� ������L# 5�Yk}���  /��6///1/C/ U/g/=�/a�/�/? �/�/D??-???�?c? u?�?�?�?�?�?�?�? @OO)OvOMO_O�O�O �O�O�O�O�O�/�/�/ __�_�Om__�_�_ �_o�_�_8oo!o3o EoWoio�o�o�o�o�o �o�o�ojAS �;_M_{��u� ���+�x�O�a��� ��������͏ߏ,�� �b�9�K�]�o����� ����ɟ����� p��Y�k�������� ůׯ$�����l�C� U���y���ؿ����ӿ  ���	�V�-�?ό�'� 9�K�yϋ�a�����.� ��d�;�M�_�q߃� ���߹�������� %�7�I��m����� �����&�������� E�W���{��������� ������X/A� ew����� �B+=��7� ew���/�/ P/'/9/K/�/o/�/�/ �/�/?�/�/�/L?#? 5?�?Y?k?�?�?�?�? �O��?�?ZO1OCO �OgOyO�O�O�O�O_ �O�OD__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo)o�?�o#OQoco �o�o�o�o�o %7�[m��� ����8��!�n� E�W�i�{�����uo�� �oǏُF��/�|�S� e�w�ğ������џ� 0���+�x�O�a��� ����䯻�ͯ߯,�� �����=�O���7� ����ɿۿ�:��#� p�G�Y�k�}Ϗϡ��� ����$�����1�C� Uߢ�yߋ���s����� ��2���-�?�Q�c� ������������� ��d�;�M���q��� ����������N ����);�#�� ���&�\3 EW�{���� /��/X///A/�/ e/w/�/_q��/�/ �/??f?=?O?�?s? �?�?�?�?�?O�?O PO'O9OKO]OoO�O�O��O�O_�O�O�O�$��$DCSS_PS�TAT ����cQQ �   t_�Z r_ (�_�_�WkP�kP�_�_ l 	cdP��P;_4oFo�)"ocUcUdovoTT�SETUP 	NcYB�&T�#�!��dOYT1SC 2i
�j`�!Cz�#�/}�eCP R-�l�� DSoz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ��.h%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� ������������ +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G��� ��}������������� ��1CUgy �������	 -?Qcu��@�����Z�D�/ */</�/`/r/�/S/�/ �/�/�/�/??�/8? J??[?�?�?a?�?�? �?�?�?O"O�?FOXO jO9O�O�O/}O�O�O oO__0_�OT_f_x_ G_�_�_�_�_�_�_�_ o,o>ooboto�oUo �o�o�o�o�o�o :L�O)��� ��� ��$��H� Z�l�;�����q���؏ ꏹ�� �2��V�h� z�I���������� _՟.�@�ǟd�v��� W�����Я������ �<�N��_�����e� ��̿޿����&����J�\�n�=ϒϤ�s���$DCSS_TC�PMAP  ������Q_ @ ~�~��~�~���~��~�~�~�	g� � ~�~�~��~�~�~�~��~�~�~�~�J~�~�~�~�~�U~�~�~�~�U~� ~�!~�"~�U#~�$~�%~�&~�U'~�(~�)~�*~�U+~�,~�-~�.~�U/~�0~�1~�2~�U3~�4~�5~�6~�U7~�8~�9~�:~�U;~�<~�=~�>~��?~�@��UIROw 2�����$��"�4�F�X�j� |������������@��0�B�T�}�� }������������� 1CUgy� ����^����� -?Qcu��� ����//)/;/ M/_/��/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�?�v/O��UIZN �2��	 ��� ��PObOtOy�KO�O�O �O�O�O�O_�O0_B_ T__x_�_�_k_�_�_ �_�_�_o,o�_Pobo to�oIo�o�o�o�o�o �o:L^-� ��i����� $�6��Z�l�~�M��� ��Ə؏�����ݏ2��D�V�O��UFRM; R������ ����ß՟����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� ���߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��ߗ����� ������'9K ]o������ ��#5GYk���x���� ��//�B/T/// x/�/e/�/�/�/�/�/ �/?,??P?b?y� �?�?I?�?�?�?OO �?:OLO'OpO�O]O�O �O�O�O�O�O�O$_6_ _Z_l_�?�_�_A_�_ �_�_�_o�_2oDoo hozoUo�o�o�o�o�o �o�o.	Rd{_ ��9����� ��<�N�)�r���_� ������ޏ��ˏ�&� �J�\�sw