��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�ASSNAME_�T   0 }$+ $'�WORD  ? L�EVEL  w$TI- OUTT� &F/�� $SETUP�JPROGRAM�JINSTALL�JY  $C�URR_O�US�ER�NUM�S�TPS_LOG_ZP N��$�T��N�  6 CO�UNT_DOWN��$ENB_PCMPWD � �DV�IN!s$C� CRE�OPARM:� T:DIAG:)��LVCHK!F�ULLM0�YX=T�CNTD��MENU�AUT�O,�FG_DS�P�RLS����$$CL(   O���!��	���	�$DCS_C�OD@���%��  W'_S � *�! V&��A91("!�0 d $VA�G M/��R�J3ICSPEZ�VW���   5?67 TOR�$�#�P� ��!LINEBUILD�"?2007�%���� FANUC���25111�7 7�� 
BEDIEN�% 0O�&T �!�J006�'  7599���"6�&K=:708;9608m;43�J7D1292�?10v�:27�?011�%=�� 9303�6�"x�2�4�38085�?I1�7�14I5J4�9�235HG"G�154�jO01:4�3653r"O00�8003:4�w�G�4�D09p�4JFG� 118G2F2�G�A36ZG(Wn�:597�O02J�098�G(W6J42�5�_02ZJ793��7(W~J50Y(W�J4�16�G(W�J7666�_02�J49}H(WnZ493_032Z�794o0�X�A1�_�`J16_�`�[�45B_03ZJ10��o�`~J2�Y�g�J1�57FO03�K29v�o03�J734bo�03Z06�_J0m4�k78�_04�;�18�o04J367�0�H�!�?�qZJ�94	h�w~J817��0�h�Q85�0�4�J13�8�w�K2H)x�wZ73�3�52Z�54�J10�:22UX��J����6J����ZJ59H��N{� ���J+����JO����J s���Z�����5��Ǩ���䯲��֟��{510�_�ZJ43ŏ_�bN{9��ȧ�J99���Ϡ�L��ȧ[7A_J�11[49�5-��:3�8��0��35J�1.�[575Z�1�[��:��1�U���RyX�0�r{1i�0�λ86���1QkL���1uk5k85~�1�k47E��`��;8�h`�J66 �������qxX����D^�J5c�C�q{9�iDX��J3<o^�Rk8��_�Z8[p���8850��1%�82���J46��>�d�ZK ������B���f������
B�J4w 
��PDonpro�$�T�΀vEG.!b#SU»!n+�/�/b#WORD �!�9t�n;0  
�1d,4 V�[t&��j1�10CB ����