A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �SBR_T   | 	$SVMTR_ID  $ROBOT_ID $GRP_NUM  $AXIS_NUM  $MTR_ID $MTR_INF_ID $SV_PARAM_ID 	$PARAM  ,$MOT_SPD_LIM    �SBR2_T   $PARAM   �  D�$$CLASS  ������       �$SBR 1 ������ T�    M-900iA/260L                aiS30/4000 160A       
H1 DSP1-S1    	P01.04    ,  	�     Pa       ���   ��    
=  
	��r9  ��9 :    D 8HB  �����         � �                  ��         3!��=����3�n%d
�                 & ���� t      �S                       �F��        E��;����	�         YB� S K     S �	� :?O�        'b��                                                                                                                                                                                                                                                                                                     �    M-900iA/260L                aiS40/4000 160A       
H2 DSP1-S2    	P01.04    ,  	�     Pa       �����   �$    
=  
8�'r9  c��9 :    D @mB ,��	`� �        y t                  �l         3�p��=������i�                   ���� U      �u                       ���S        
����3b���         �B� � H     � �� :?=�          �	                                                                                                                                   3                                                                                                                                                                  �    M-900iA/260L                aiS40/4000 160A       
H3 DSP1-S3    	P01.04    ,  	�     Pa       �����   ��    
=  
8��r9  c��9 :    D @mB ,��@� �        y 8                  �k         8� ��8/����V�
�                   ���� 3      ��                       ���J        ��U�����        �B� � H     � �� :?=�          �	                                                                                                                                   	�                                                                                                                                                                  �    M-900iA/260L                aiS12/4000 40A        
H4 DSP1-S4    	P01.04    ,  	�     Pc        �q��   2�$    {  
8�(r9  ~�k0�        � (H�  ���	`��/        �                  �                                                     / ���� ]      ��                       B�W         ?��
��h��         �a  6     �� :?�          y/                                                                                                                                  f                                                                                                                                                                  �    M-900iA/260L                aiS12/4000 40A        
H5 DSP1-S5    	P01.04    ,  	�     Pc        �q��   2�$    {  
8�'r9  ~�k0�        � (H�  ���	`��        � �                  �                                                     5 ���� a      ��                       L��         ��
+����\q        <a  6     �� :?�          y/                                                                                                                                  f                                                                                                                                                                  F    M-900iA/260L                aiS12/4000 40A        
H6 DSP1-S6    	P01.04    ,  	�     Pc        �q��   2�H    
=  
8�Nr9  ~�k0�        � (H�  ���	`��:       � �                  �                                                     " ���� `      �%                       �	N         ��X	��{�         �a  6     �� :?�          y/                                                                                                                                  f                                                                                                                                                                  m����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$SBR2 1������ T0 �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������