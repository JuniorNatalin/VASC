A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �SBR_T   | 	$SVMTR_ID  $ROBOT_ID $GRP_NUM  $AXIS_NUM  $MTR_ID $MTR_INF_ID $SV_PARAM_ID 	$PARAM  ,$MOT_SPD_LIM  ��SBR2_T   $PARAM   � ��$$CLASS  ������       �$SBR 1 ������ T�    R-2000iB/210F               ACaiSR30/3000 80A     
H1 DSP1-S1    	P01.05    ,  	�     PaR�      ����   �    
=  
#�,r9  ~��%�9      8 l�  ����� %        �(       ��      �k   �/  3!���=�����=��vG��          &��S  ���� m      �                       ���Z        	��y	��y��j�         �c9	`B 0     � �� :?p�   @  'bx�                                                                                                                                  3                                                            Z                 3!���=����e��3@���=���� 
�'�!                                          ,    R-2000iB/210F               ACaiSR30/3000 80A     
H2 DSP1-S2    	P01.05    ,  	�     PaR�      ����   �@    
=  
8�Dr9  ~��%�9      8 l�  ����� h        � �               ��   �� 3�f��<����wD��7�D          &��#  ���� O      �S                       ����        ��2��2
��(�         �c9	`B 0     � �� :?p�   @    x�                                                                                                                                  3                                                            Z                 3E���=����N	5�5k
}��;w�/��
�
k'�:                                              R-2000iB/210F               ACaiSR30/3000 80A     
H3 DSP1-S3    	P01.05    ,  	�     PaR�       ����   �\    
=  
3�cr9  ~��%�9      8 l� �p��� h        � y       /�/�       ��         3����<����F�4���D          &�      ���� 6      �v                       ���K        	��	��9��S�         �c9	`B 0     � �� :?p�   @    x�                                                                                                                                  3                                                            Z                                                                                                   �    R-2000iB/210F               ACa12/4000iS 40A      
H4 DSP1-S4    	P01.05    ,  	�     Paz       �q��   2�m    
=  
8�pr9  ~�k0�        � (H�  �������        � �       @@      �                                                      ���� ;      ��                       ���0         ]���VP��        ��       �� :?�          y/                                                                                                                                  f                                                                                                                                                                  �    R-2000iB/210F               ACa12/4000iS 40A      
H5 DSP1-S5    	P01.05    ,  	�     Paz       �q��   2��    
=  
8��r9  ~�k0�        � (H�  ������
�        �       >�>�      �                                                      ���� :      ��                       ���         N�P���9        ��       �� :?�          y/                                                                                                                                  f                                                                                                                                                                  �    R-2000iB/210F               ACa12/4000iS 40A      
H6 DSP1-S6    	P01.05    ,  	�     Paz       �q��   2�     
=  
8�$r9  ~�k0�        � (H�  �������        � �       LL      �                                                     * ���� 9      ��                       ��         ��<��
��U�       .�       �� :?�          y/                                                                                                                                  f                                                                                                                                                                  M����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$SBR2 1������ T0 �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������