A��*SYSTEM*   V8.2306       4/24/2014 A5  *SYSTEM*  ��AAVM_WRK_T  � $EXPOSURE  $CAMCLBDATE $PS_TRGVT   $TRGVT  $TRGHZ  $TRGDIST  $TRGW  $TRGP  $TRGR  $LENS_CENT_X  $LENS_CENT_Y  $DISTORT   $CMP_GC_P  $UTNUM  $PRE_MAST_CT   	$PRE_GRV_MST  $NEW_MAST_CT   	$NEW_GRV_MST  $STAT_RUN  $RES_ERR  $VTCP_ERR   $TRGT_ERR   $RES_ERR2  $VTCP_ERR2   $RSM_MAST_CT   	$STAT_START  $STAT_END  $STAT_ORGBK  $STAT_RSMBK  $STAT_ORGRES  $STAT_UPDT  �ABSPOS_GRP_T   $PARAM   
x�ALRM_RECOV_T    $ALMRECOVENB   $ALMRECOVON   �ALMDG_T  0 $DEBUG1  $DEBUG2  $DEBUG3  $CONT_TYPE  �ALM_IF_T  D $ENABLE  $LAST_ALM d$LAST_UALM d$KALM_MAX  $LDEBUG   
 ��APCOUPLED_T  $ $APP_PROCES0  $APP_PROCES1   ��APCUREQ_T  � $SOFTPART_ID  $TOTAL_EQ  $CUR_EQNO  $PS_SPI_INDE   $SPI_INDEX  $SCREEN_NAME $APP_SIGN $APP_PROCES0  $APP_PROCES1  $TOPK_FILE 	$THKY_FILE 	$PANE_EQNO   	$DUMMY12  $DUMMY13  $DUMMY14  ��ARG_STR_T  � $TITLE $ITEM1 $ITEM2 $ITEM3 $ITEM4 $ITEM5 $ITEM6 $ITEM7 $ITEM8 $ITEM9 $ITEM10 $ITEM11 $ITEM12 $ITEM13 $ITEM14 $ITEM15 $ITEM16 $ITEM17 $ITEM18 $ITEM19 $ITEM20 
��ASBN_CFG_T  8 $CNV_JNT_POS  $DATA_CMNTS  $FLAGS   $POS_CHECK  �AT_CELLSETUP 	 P $HOME_IO_PRG %$HOME_MACRO %$REPR_MACRO %$PRODRUN_SPD  $PRODRSM_SPD   �AUTOBACKUP_T 
 $ENABLE  $DEVICE $TIME   $DI_IDX  $STARTUP_BCK  $INTERVAL  $DISP_UNIT  $BCK_DO_IDX  $ERR_DO_IDX  $FR_FREE  $IN_PROGRESS  $REQ_BACKUP  $PRC_WAIT  $AUTO_BACKUP  $POFF_COUNT  $DEL_COUNT  $LOG_IDX  $DEL_TIME ? $DEL_FILE ?� $PROC_FILE ���MOTOR_COUNTE  0 $REM_COUNTS   	$REM_REV   	$BIL_REV   	,�AXIS_COUNTER   $ODOMETER $NON_CMD ��AXIS_METER_T    $ODOMETER   	$NON_CMD   	��AXSCRDCFG_T  d $CARD_EXIST  $FSSB_TYPE  $CHKBD_SEL  $DIAG_REG   $SLOT_NUM  $SLOT_PREV  $DEBUG   8�BACK_EDIT_T  � $PROGRAM %$SRC_NAME %$EPT_IDX  $OPEN_ID  $DELETE_OK  $USED_TP_CRT  $BACKUP_NAME %$PS_REPLACIN   $REPLACING  $BCK_COMMENT $D_REPLACING  $SEL_PROGRAM %$DUMMY12  $DUMMY13  ��BLAL_OUT_T  , $DO_INDEX  $PS_BATALM_O   $BATALM_OR  �CFCFG_T  X $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $COMP_SWITCH  $MAX_NSETS  �CF_PARAMGP_T  � 
$WARNMESSENB  $CHKJNTLIM  $CNSTNT_CORN  $TIMEFLTRENB  $TRATIO_TB   $ACCTIME_TB1   $ACCTIME_TB2   $ORIENT_TYPE  $DEBUG  $RTSPD_SF  ��CHG_PRI_T   $TASK_ID  $PRIORITY  ��CHKPOS_T  x $CONT_FLAG  $POS_HDR  $JPOS1  $JPOS2  $JPOS3  $JPOS4  $JPOS5  $JPOS6  $JPOS7  $JPOS8  $JPOS9   ��COCFG_T  < $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $ENABLED  �CO_MORGRP_T  t $FLEN  $ANGLE  $TBA_MAG  $TBA_MAG_PRE  $TBA_MAG_MAX  $TBA_MAGAXS   	$TBA_CURAXS   	$TBA_PRVAXS   	��CO_PARAMGP_T  � $OPT_TIME  $OPT_ACC  $JACC_RRATIO  $CACC_RRATIO  $JTIME_RATIO  $CTIME_RATIO  $JVARDMAX  $CVARDMAX  $WARNMESSENB  $DEBUG  $TBA_MGN  M��CP_RSMOFST_T  @ $RO_ENABLE  $RO_MAX_ITP  $RO_NOM_DIST  $RO_NOM_SPD   ��CPCFG_T  � $GROUP_MASK  $CP_DEBUG  $CP_ENABLE  $COMP_SWITCH  $EXTRA_INT   $EXTRA_FLT   
$TF_MODE  $MD3ITPTOL  $RESUME_OFST $CP_HSTART  $T1_HSTART  $TEST   $COMP_SW2  $COMP_SW3  $COMP_SW4  ��CPDBGDEF_T  d $OUTPUT  $FILENAME )$GROUP_MASK  $DEBUGMASK  $MAXDATA  $COUNT  $TAIL  $BUFEXIST  `�CPDBG_T  � $OUTPUT  $CPIDEBUG $CPPDEBUG $MIDEBUG $MPDEBUG $MGDEBUG $MFDEBUG $SIMQSTOP  $KEEP  $PATH )$EXTRA1  $EXTRA2  ��CP_L64FIX_T  � $ENABLE  $DEC_A   $DEC_V   $DEC_CIF   $DEC_PCHO   $ADD_A   $ADD_V   $ADD_CIF   $ADD_PCHO   $DEBUG_SIM  $SIM_ADDRESS  $SIM_VAR_TYP  $SIM_AXIS  $EXTRA1  $EXTRA2  $EXTRA3  ��CP_MCRGRP_T  4 $RSM_JBF_PCT  $RSM_DEC_PCT  $RSM_OFS_PCT   D�CP_MORGRP_T  � $CHNS_EMPTY  $GTF_EMPTY  $CHK_T1_SPD  $T1_FPSPD  $T1_TCPSPD  $SPEED  $T1SPDLIM  $SPEEDTOL  $JNT_VEL   	$JNT_ACC   	$JNT_JRK   	$SEGFRACTION  $RSTRT_LINE  $RSTRT_PVF  H�CP_TESTDEF_T    $ENABLE_TEST  $NUM_LINES  X�CP_PARAMGP_T  D )$WARNMESSENB  $DEBUG  $ENB  $NUM_CHN  $NUM_JBFSET  $NUM_JBF  $EXT_NUM_JBF  $JBF_SIZE  $EXT_JBF_SIZ  $NUM_TF  $TF_SIZE  $EXT_TF_SIZE  $NUM_RSINFO  $JNT_VEL_LIM   	$JNT_ACC_LIM   	$JNT_JRK_LIM   	$T1SEGFL_SF  $T1GTFL_SF  $CRCMP_SWITC  $ACCLIM_SF  $JRKLIM_SF  $PSPD_SWITCH  $MAX_PSPD  $MIN_PSPD  $PSPDACC_SF  $PSPDJRK_SF  $CDCOMP_SW  $CDACC_SF  $CDJRK_SF  $CDDELTATOL  $CDDISTSF  $CDANGTOL  $CDDEVTOL  $CHKJNTLIM  $FDANG_TOL  $FDLIN_TOL  $JNTJBF_ENB  $COMP_SW  $EXTRA_INT   $EXTRA_FLT   $CP_TEST <�CP_T1_MODE_T ! � 	$ENABLE  $COMP_SWITCH  $MARGIN  $TIME_FACTOR  $SPD_LIMIT  $SLEW_RATE  $MIN_TFLEN  $EXTRA_INT   $EXTRA_FLT    l�CRCFG_T "� $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $PGDEBUG  $CR_ENHANCED  $LGORN_ENBL  $BLEND_ENB  $MAX_ARC_ANG  $RSM_RSPD_LM  $LGORN_METH  $LGORN_DBG  $LGORN_RAD  $LGORN_AZ_SP  $LGORN_ELTOL  $ROTSPDFCTR  $MAX_FP_SPD  $SMCRC_RADI  $SMCRC_RADO  $SMCRC_ARC  $ARCANGLIM  $MAXORNTCHG  $MAXSGRATIO  $CHKBMP  $RSM_TYP  $CHK_MSK  $AES_SINGTOL  ��CRI_CFG_T #  $CRI_SW  �CSXC_PARAM_T $ x 	$NAME $ATTR  $NUM_CHANNEL  $IMG_HEIGHT  $IMG_WIDTH  $VT_SPACING  $DEF_ASPECT  $MIN_EXPO  $MAX_EXPO  �CUSTOMMENU_T % $ $TITLE $PROG_NAME %$OPTION  �CZ_CDCFG_T & x $ENABLE   $CD_ENABLE  $NO_HEADER  $COMP_SWITCH  $WARNMESSENB  $EXTRA_INT   $EXTRA_FLT   $CHK_SPD_SF  ��DBPXWORK_T '  $SKP_DEL   U��DBTB_CTRL_T ( � $ACRT_MODE  $MINDT_ADJ  $DELAY_CALL  $DELAY_DO  $DELAY_PLS  $RESERVED1  $RESERVED2  $RESERVED3  $NUM_IO  $DUMMY9  $DUMMY10  ��DB_DBG_T )  $DBG_PRM   
��DPOS_DAT_T *  $X  $Y  $Z  t�LDPOS_DAT_T +  $X  $Y  $Z  0�PD_T ,  $X  $Y  $Z  ��PC_T -  $X  $Y  $Z  x�PENETRATE_T .  $X  $Y  $Z  @�DB_RECORD_T /H $CPOS *$LPOS +$DPOS_DST  $LDPOS_DST  $LINE_NUM  $ONCE_DC  $CROSS  $TASK_ID  $ENABLED_TIM  $TRIGGER_TIM  $PAUSED_TIME  $RETURNED_TI  $MMR_STATUS $CRE_NEWMON  $SIGNAL_ACT  $LAST_ACT  $PD ,$PC -$PN_AT .$PD2  $PC2  $PT  $PD_DOT_PC  $LINE_DST  $P_NUM  $GO_AWAY  $MOTION_COMP  �DCSS_DEVICE_ 0 P $TYPE  $RBT_NUM  $SPI_IDX  $SPO_IDX  $SPI_BYTE  $SPO_BYTE  $STO  �DCSS_LS_T 1 H $STOOUT_IDX  $STOFB_IDX  $STOFB_CH  $FENCE_TYPE  $FENCE_IDX  �DCSS_PARAM_T 2 H $DOCHK_ENB  $PMCS_ENB  $LS_STOP  $LS_FENCE  $HOTSWP_TIME   ��DCSS_ELEM_T 3 T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    	t�DCSS_RBT_T 4 � $MDL_ELEM 23 
$ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$FB_TOL   	$RBT_TYPE  ��DCS_CFG_T 5� $DISP_MENU  $LOG_ENB  $LOG_LEN  $LOG_FILE $LOG_ID  $LOG_IDMAX  $LOG_DELAY  $LOG_WRT  $LOG_INTVL  $LOG_EVENT  $TEST_PARAM1  $TEST_PARAM2  $CHK_J_TOL  $CHK_C_TOL  $SAFE_SPD  $SAFE_SPD_SV  $EXCLUDE   $SPD_ONLY   $SYS_PARAM  $PROTECT  $HI_VRC  $APPLY_WARN  $HIDE_MENU  $HI_VRC_MLT   $VRFY_ALL  $HI_MATE  $IOC_PROT  $IOC_CRC1  $IOC_CRC2  $OPI_VRC  �DCS_CRC_OUT_ 6  $START_GRP    h�DCS_SGN_T 7 � 
$CURR_SIGNAT  $CURR_DATE $PREV_SIGNAT  $PREV_DATE $ANNUNC_TYP  $ANNUNC_IDX  $CUR_TIME   $LATCH_TIME   $CUR_CRC   $LATCH_CRC    	��DEFLOGIC_T 8 @ $FUNC_TITLE 	$TOTAL_NUM  $DUMMY2  $DUMMY3  $DUMMY4  ��DEMO_INIT_T 9 L $DEMO_ENB  $DEMO_AU  $DEMO_DAYS  $LOAD_NUM  $DUMMY4  $DUMMY5  X�EFF_AXIS_T :  $NUM  $COEFF  ��ADJ_RTRQ_T ; D $COR_TRQ   $COR_TEMP   $EFF_AXIS 2: $LIMIT  $ADJ_NUM  ��AMP_COEF_T < 0 $COEF_A   	$COEF_C  $MASK  $DUAL_MASK  �CTRL_CAB_T = @ $TRANS_A  $IDLE_PWR  $AMP_COEFB  $SV_NUM  $SV_AMP 2< �DIAG_GRP_T >8 *$VAL_SET  $TACC   	$TACC_LIM1   	$TACC_LIM2   	$RRATE_LOAD   	$VER $ANSWER  $RCC_ANS  $ADJ_RTRQ 2; $ADJ_OHTRQ   	$COPPER   	$IRON   	$BRK_PWR   	$CABLE_ACT   $CABLE_BASE   	$CABLE_LENG   	$CAB_NUM  $CTRL_CAB 2= $TRQCNS   	$TRQDWN   	$MSBAS   	$MAXTRQ   	$RRATE   	$LIFECALC   	$L10   	$N0   	$T0   	$CUR_L10   	$TCP_TYPE  $CUR_TCP $MOTN_STYLE  $FLAG  $CUR_OVC   	$CUR_HEAT   	$SUPPORT_TYP   	$ALL_SUPPORT  $CUR_TCP_X  $CUR_TCP_Y  $CUR_TCP_Z  $CUR_TCP_W  $CUR_TCP_P  $CUR_TCP_R  	��DICT_CFG_T ? ` $CACHE_ENB  $CACHE_SIZE  $CURR_ONLY  $LANG_SUFFIX $LOCALE  $DUMMY5  $DUMMY6   	(�DMSW_CFG_T @ 8 $KEYIMAGE  $TMS_DSB  $TMS_STAT  $TMS_INPUT   	��DOCVIEWER_T A  $DBGLVL  $CURFILE ?� 		��DPM_CFG_T B x 
$ENABLE  $DPM_INLINE  $GRP_MSK  $BEF_JBF  $DELAY  $ORI_CTL  $CUR_SCH  $MAX_SCH  $COMP_SW  $DEBUG  (�OFS_CHN_T C � $ENABLE  $OTF_DI_IDX  $CHN_TYP  $RAMP_GAIN  $SCAN_RATE  $INI_OFS  $REM_OFS  $APP_OFS  $IN_TICK  $OU_TICK  $ID  $STAT  $MAX_LIM  $MIN_LIM  $MAX_INC  $MIN_INC  $A1  $A2    �AI_CHN_T D  $P_GAIN  $D_GAIN  $I_GAIN  $STR_CNT  $REF_CNT  $AVE_CNT  $FBK_MODE  $REF_VAL  $RAW_FBK  $CAL_FBK  $PORT_NUM  $CAL_DONE  $SLOPE  $INTERCEPT  $CUR_TICK  $LEAD_DIS  $BUF_SIZE  $BUF_CNT  $T_ADJ  $MIN_VAL  $MAX_VAL  	p�BI_CHN_T E D $DI_IDX1  $DI_IDX2  $BUMP_OFS  $BUMP_RATE  $BUMP_GAIN  ��GI_CHN_T F  $DI_IDX  $SCALE  ��DPM_GRP_T G � $OFS_TYPE  $OFS_FRAM  $LAST_DPM  $OFS_ACCU  $OFS_ABS  $OFS_CARRY  $CTL_RATE  $INT_LINE  $OFS_LINE  $DAT_RDY  $OFS_STAT  $SND_TYPE  $TRK_MODE  $SYNC_DI  $OFS 2C 	$AI_CH 2D 	$BI_CH 2E 	$GI_CH 2F 	��DPM_SCH_T H 0 $GRP_MSK  $COMMENT $DPM_ON  $GRP 2G L�DPM_IN_T I 8 $LINE_NUM  $DELAY  $OFS_X  $OFS_Y  $OFS_Z  T�DRC_CFG_T J D $HOST1 !$HOST2 !$HOST3 !$HOST4 !$HOST5 !$EMAIL_ENABL  �DSBL_FAULT_T K  $ENABLE  $MAX_COUNT  ��DTREC_T L, $DTREC_ENB  $SAMPLE_ITP  $BUF_SIZE  $FILE_SIZE  $DEVICE_NAM $SUBBUF_SIZ  $SPC_FILE  $DTREC_ON  $DTSAV_ON  $FILE_ACCESS  $PC_ACCESS  $SYSTIME   P$DTSAV_ENB  $ORDER  $DSB_BUFSIZ  $ENB_BUFSIZ  $OTTASK_MOD  $DP_ALM_ID  $DP_ALM_GRP  $DP_ALM_AXS  $DEF_MAXBUF  |�DYN_BRK_T M 0 $DI_IDX  $DO_IDX  $BRK_MSK  $FLTR_IF  ��ENC_STAT_T N� $ENC_COUNT  $ENC_ROS_TIK  $ENC_RATE  $ENC_AVERAGE  $ENC_ENABLE  $ENC_DSPSTAT  $ENC_SPCSTAT  $ENC_SIM_ON  $ENC_SIM_SPD  $ENC_VALUE  $ENC_HEAD  $ENC_MULTIPL  $ENC_STOPPED   $ENC_THRESH  $ENC_EXISTS  $ENC_HSDI  $ENC_ABSCNT  $INCTRAVDIST  $INCTRAVCNTS  $INCTRAV_DO  $CONVSPD_GO  $INCTRAVRES  $ENC_BUFFER   d$ENC_ATR_AXS  $SC_GRP_NUM  $ENC_COMERCT  $ENC_FBCMPCT  �ENETMODE_T O 8 $FULL_DUPLEX  $SPEED  $ACD_ENABLE  $THROTTLE  ��ER_NOAUTO_T P D $NOAUTO_ENB  $NOAUTO_NUM  $PS_NOAUTO_C   $NOAUTO_CODE    x�ER_NOALM_T QH *$NOALMENBLE  $NOALM_NUM  $ER_CODE1  $ER_CODE2  $ER_CODE3  $ER_CODE4  $ER_CODE5  $ER_CODE6  $ER_CODE7  $ER_CODE8  $ER_CODE9  $ER_CODE10  $ER_CODE11  $ER_CODE12  $ER_CODE13  $ER_CODE14  $ER_CODE15  $ER_CODE16  $ER_CODE17  $ER_CODE18  $ER_CODE19  $ER_CODE20  $ER_CODE21  $ER_CODE22  $ER_CODE23  $ER_CODE24  $ER_CODE25  $ER_CODE26  $ER_CODE27  $ER_CODE28  $ER_CODE29  $ER_CODE30  $ER_CODE31  $ER_CODE32  $ER_CODE33  $ER_CODE34  $ER_CODE35  $ER_CODE36  $ER_CODE37  $ER_CODE38  $ER_CODE39  $ER_CODE40   ��ER_OUTPUT_T R � $OUT_NUM  $IN_NUM  $PLCWARN  $GRP_STR  $ERROR_NUM  $FAC_NUM  $SEV_NUM  $PARM1_NUM  $PARM2_NUM  $DUMMY9  $DUMMY10  $DUMMY11   �EXT_SET_T S < $ENABLE  $DI_TYPE  $DI_NUM  $DO_TYPE  $DO_NUM  ��FDR_GRP_T TT $VEL_MOD   	$VEL_CNT   	$REM_LIFE2   	$OVM_RATE   	$OVA_RATE   	$TROV_RATE   	$DTAV_RATE   	$DTMX_RATE   	$DTMIN_RATE   	$MOT_RATE   	$DIAG_INDX_R   
$DIAG_INDX_I   $DG_MAXT   	$DG_T0   	$RATED_TRQ   	$DRIVE_TYPE   	$GEAR_RATIO2   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$Z_MCMD   	��FEATURE_T U , $NAM ? $MOD ? $VER ? $MEC ?  �FILECOMP_T V  $TPP  $VARIABLE  ��FILE_SETUP2_ W 4 $FILE_TDC_SC  $FILE_TV_SEC  $FILE_TVC_SC   x�FILE_BACK_T X T $FILE_NAME )$PROG_NAME %$FUNC_CODE  $MODIFIER  $COMMENT %$FUNC_PTR   	��FMR2_GRP_T Y $VEL_ROT  $VEL_LIN  $VEL_MOD   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$TROV_MAX   	$T_LIFE_0  $RATED_TRQ   	$LIMIT_FUNC  $ACC_LMT   	$DRIVE_TYPE   	$GEAR_RATIO2   	$DGCLFR   	$DGDYFR   	$DGLDEC   	$DG5T0   	$DG_MAXT   	$DG_T0   		��FMR_CFG_T Z  $TROV_MAX   T�FSSB_CFG_T [ P $FSSB_LINE   $EX_FSSBLINE   $FSSB1_AXES  $FSSB3_AXES  $FSSB5_AXES  �GRAVC_GRP_T \ � 
$MODE_SW  $SPCONS   	$DEBUG1  $DEBUG2   	$GRV_STATUS  $BKUP_NO116   	$POFF_NO116   	$GRVCMP_SW  $GRVMST_LOOP  $MST_SMT_LEN   H�MOTYPE_E ]       �TERMTYPE_E ^      d�ORIENT_E _       �SM_PROFILE_E `      �TA_PROFILE_E a       �UPR_T b� -$MOTYPE ]$TERMTYPE ^$SEGTERMTYPE ^$DECELTOL  $USE_CONFIG  $USE_TURNS  $ORIENT_TYPE _$UFRAME $UTOOL $SPEED  $ROTSPEED  $CONTAXISVEL  $CNSTNT_PATH  $CNSTNTPTHJT  $SEG_TIME  $USE_CARTACC  $USEMAXACCEL  $USERELACCEL  $USETIMESHFT   $USE_PATHACC  $USE_SHORTMO  $SM_PROFILE  `$TA_PROFILE  a$ACCEL_OVRD  $TIME_SHIFT  $ACCU_NUM   $PAYLOAD  $DYN_I_COMP  $PATHRES_ENB  $RESERVE1   $CNT_SHORTMO  $EXT_SPEED  $CNT_ACCEL1  $CNT_ACCEL2  $CRCCOMPENB  $ASYMFLTRENB  $USE_WJTURNS  $EXT_INDEP  $CARTFLTRENB  $CNT_SPEEDUP  $CNT_DYN_ACC  $MAX_SPEED  $USERELPSPD  $PSPD_OVRD  $ORNT_MROT  ��GRSMT_GRP_T c  $GRV_SW  $GRV_PARAM  l�HOST_CFG_T d � $COMMENT $PROTOCOL 	$PORT $OPER  $STATE  $MODE $REMOTE $REPERRS  $TIMEOUT  $PATH e$STRT_PATH e$STRT_REMOTE $USERNAME e$PWRD_TIMOUT  $SERVER_PORT  $USE_VIS_PRT  ��HOSTENT_T e 4 $H_NAME !$H_ADDRTYPE  $H_LENGTH  $H_ADDR !T�ERR_MASK_T f H $SSC_MASK1  $SSC_MASK2  $SSC_MASK3  $SSC_MASK4  $SEV_MASK  h�HSCD_MNG_T g $COLL_MODE  $THRESHOLD  $DO_ERR  $DO_ENABLE  $MACRO_REG  $STND_CD  $AUTO_RESET  $UPD_GROUPS  $PARAM_VERID 	$PARAM119   	$PARAM120   	$PARAM121   	$PARAM122   	$PARAM123   	$PARAM124   	$PARAM125   	$ACT_RATIO  $SAVED119   	$SAVED120   	��HSCD_GRP_T h $ $COL_DET_OFF  $HSCD_PRM_ID  T�HTTP_AUTH_T i ( $OBJECT !$NAME $TYPE  $LEVEL  �HTTP_T j � $ENABLE  $ENAB_DIAGTP  $ENAB_SPART  $DBGLVL  $KRL_TIMOUT  $HITCOUNT  $BG_COLOR $ENAB_TEMPL  $TEMPLATE $COMMENT $RSS_INUM  �HWR_CONFIG_T k H $MAINCPU  $VISIONCPU  $SPARE1  $SPARE2  $SPARE3  $SPARE4  `�IBGN_CFG_T l $CMP_WAIT  $MAX_PNUM1  $MAX_PNUM2  $FWD_TOL_LOC  $FWD_TOL_ORT  $FWD_TOL_EXT  $FWD_TOL_ANG  $BWD_TOL_LOC  $BWD_TOL_ORT  $BWD_TOL_EXT  $BWD_TOL_ANG  $BWD_RTN_SPD  $UF_DATA  $DBG_MASK  $TEMP_MGN  $LIN_N_CNST  $END_TOL_LOC  $STATUS  $RECDAT_SEND  8�IBGN_ERRIO_T m @ $REC_IO_TYP  $REC_IO_NUM  $EXE_IO_TYP  $EXE_IO_NUM   |�IBGN_EXEC_T n ( $SCHEDULE   $FILE_P   $BWD_FLG    <�IBGN_FIL_T o @ $EXE_MD  $EXE_OPN  $EXE_BACK  $REC_TRANS  $REC_ACC  d�IBGN_FTP_T px $FTP_CTAG  $AUTO_TRANS  $IGNR_COMER  $FTP_STAG  $SM_STAG  $SM_CTAG  $SM_SPORT  $SM_CPORT  $N_PCSOFT 	$N_RECFL1 	$N_RECFL2 	$N_RECFL3 	$N_EXEFIL $N_FLEXT1 $N_CONDFL 	$N_FLEXT2 $N_SPTXT1 $N_SPTXT2 	$SEQ_VAR  $SNS_NUM  $SNS_CNST  $FOLDER $RECS_PRG %$RECS_TMO  $RECE_PRG %$RECE_TMO  $SM_DBG  $AUTO_START  $RESERVE  ��IOLNK_T q 8 $RACK  $SLOT  $INPUT_N  $OUTPUT_N  $OPTION  ��IOSLAVE_T r  $INPUT_N  $OUTPUT_N  \�IO_DEF_ASG_T s T $LOG_TYPE  $LOG_NO  $NUM_PORTS  $RACK  $SLOT  $PHY_TYPE  $PHY_NO   H�IO_UOP_CFG_T t ` $UOP_TYPE  $IN_RACK  $IN_SLOT  $IN_STRTPT  $OUT_RACK  $OUT_SLOT  $OUT_STRTPT   ��UJR_GRP_T u � $FINE_OVRD  $JOGFRAME $FINE_DIST  $J7_GROUP  $J8_GROUP  $J7_AXIS  $J8_AXIS  $J7_LABEL $J8_LABEL $J7_GRAPHIC Q$J8_GRAPHIC Q$DSB_J7J8  $DSBL_KEY   �KAREL_CFG_T v 0 $CONV_ENABLE  $CONV_CTRL  $CONV_FLAGS  8�LGCFG_T w � $ENABLE  $OUT_SW  $LG_SIZE  $EV_SIZE  $MR_SIZE  $SG_SIZE  $FD_SIZE  $MI_SIZE  $ER_SIZE  $MP_SIZE  $MG_SIZE  $PE_SIZE  $LG_MODE  $EV_MODE  $MR_MODE  $SG_MODE  $FD_MODE  $PE_MODE  $EX_RSCH_FIL $COMP_SW   �LN_DISP_T x ` $HIDE_LINE_N  $DISP_MENU  $HIDE_PARLN  $HIDE_DAULN  $HEAD_PARENT $HEAD_DAUGHT  ��LOGBOOK_T yt B$NUM_ER_ITM  $NUM_ER_TYP  $NUM_REC_TYP  $NUM_SCRN_FL  $NUM_DIO  $SRAM_MARGIN  $DRAM_MARGIN  $OPTION  $LOG_ER  $LOG_ENT  $LOG_SEL  $LOG_WIN  $LOG_MENU  $LOG_JGMU  $LOG_MNCHG  $LOG_FNKEY  $LOG_JGKY  $LOG_PRGKEY  $LOG_UFKY  $LOG_OVRKY  $LOG_FWDKY  $LOG_HLDKY  $LOG_STPKY  $LOG_PRVKY  $LOG_ENTKY  $LOG_ITMKY  $LOG_RSTKY  $LOG_HELPKY  $LOG_OVR  $LOG_CRD  $LOG_STEP  $LOG_GRP  $LOG_SGRP  $LOG_UF  $LOG_UT  $LOG_FILE  $LOG_WTRLS  $LOG_PGCHG  $LOG_SETPOS  $LOG_TPKY  $LOG_DIO  $LOG_STMD  $LOG_FOCUS  $LOG_PRGEXE  $LOG_TUIKEY  $IMG_ENT  $IMG_SEL  $IMG_WIN  $IMG_FNKY  $SAVE_FILE 	$SCRN_FL  $SCRN_NO_ENT  $ANALOG_TOL  $AVAILABLE  $CLEAR_ENB  $DCS_HI1  $DCS_HI2  $DCS_HO1  $DCS_HO2  $DCS_SI  $DCS_SO1  $DCS_SO2  $DCS_OPTION  $IGNR_SAVE  $FNKEY_FLTR  $DCS_DEV  ��LOG_BUFF_T z 0 $TITLE $SIZE  $MEM_TYPE  $VISIBLE    D�LOG_STAT_T { 0 $TICK  $SPD  $POS1  $POS2  $POS3   t�LOG_DCS_T | � $ENABLE  $SPD_TOL  $OUTPUT_TYP  $OUTPUT_IDX  $GRP_NUM  $POS_TYP  $AXIS_NUM  $STOP_READY  $STOP {$ESTOP {$CSTOP {$ESTOP_DIFF {$CSTOP_DIFF { |�LOG_DIO_T } L $RACK  $SLOT  $MOD_TYPE  $PORT_TYPE  $START_PORT  $END_PORT  ��LOG_SCRN_FL_ ~  $SP_ID  $SCRN_ID   �MCSP_T  � $CLDPOP_ENB  $TRQLIM_ENB  $JOGLIM_ENB  $CLDPOP_FLG  $CLDGRP_FLG  $CLDREL_FLG  $CLR_CLDFLG  $JOGLIM_FLG  $ORGJOG_OVR  $COMP_SW  $RESERVE1  $RESERVE2  $RESERVE3  t�MCSP_GRP_T � � 	$JOGLIM_OVR  $TRQLIM_FLG  $SV_PTLIM   	$ORG_PTLIM   	$ORG_RCLMC   	$RESERVE1  $RESERVE2  $RESERVE3   	$RESERVE4   	 ��MISC_GRP_T � d $HPD_TRQ   	$DSTB_MAX   	$DSTB_MIN   	$DSTB_MAXENB   	$DSTB_MINENB   	$DSTB_EXCESS   ��MISC_MSTR_T �  $HPD_ENB   @�MISC_SCD_T � H $DSTB_MAX_A   	$DSTB_MIN_A   	$DSTB_MAXENB   	$DSTB_MINENB   	 �MKCFG_T � \ $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $MO_CONFLICT  $MO_REQUIRED  $DEBUG  0�MLTARM_CFG_T �  $NUM_ARMS  $GROUP   �MLT_GRP_DO_T � � $TP_ENABLE  $JOG_GROUP  $LOCKED_ARM  $CRNT_TYPE  $CRNT_INDX  $PRG_ROUT_P  $JOG_ROUT_P  $PRG_DO_TYPE   $PRG_DO_INDX   $JOG_DO_TYPE   $JOG_DO_INDX    ��MNDSP_MST_T � ` $DISP_ENABLE  $DISP_EDCMD  $DISP_INAUTO  $DISP_RSMDIS  $DISP_IS_ON  $MODE_GRP    �MNDSPPSTL_T � 4 $LOCTOL  $ORIENTTOL  $EXTTOL  $ANGTOL   	 ��MODAQ_CFG_T � d $ON_LINE  $MF_FLAG  $MI_FLAG  $GRP_NUM  $STARTLOG  $ENDLOG  $LN_MASK  $SUPPORT   ��FX_TRIGGER_T � � 	$START_MODEL  $START_STEP  $START_PROG %$STOP_MODEL  $STOP_STEP  $STOP_PROG %$AXES  $DATA_TYPE  $DATETIME   ��MODEM_INF_T � t $MDM_INIT )$MDM_INIT1 )$MDM_RESET )$MDM_HANGUP )$MDM_DIAL )$MDM_ANSWER )$MDM_STATUS )$MDM_IDENT )��MOR_GRP_SV_T �  $CUR_SV_ANG   	 ��ARMLOAD_T �  $ARMLOAD   ��ARMLOAD_P_T �  $ARMLOAD_P     ��MRR2_GRP_T �� $ARM_PARAM   d$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$RLIBSW01  $RLIBSW02  $ABC_FLAG  $MD_J2SECT   $MD_J3SECT   
$MD_J1SPCONS   P$MD_J2SPCONS   P$MD_J3SPCONS   P$MD_CUR_K   $MD_CUR_J2  $MD_CUR_J3  $SV_OFF_TIM2   	$CSKPLIM_ENB  $CSKPLIM_LIN  $CSKPLIM_JNT   	$QSKPLIM_ENB  $QSKPLIM_LIN  $QSKPLIM_JNT   	$EXT_AZIM   $EXT_ELEV   $SERVOCMPTOL   	$ARMLOAD 1� $ARMLOAD_X 1� $ARMLOAD_Y 1� $ARMLOAD_Z 1� ��INTERACT_T �  $INTERACTION   	t�INTRAC_N_T �  $INTRAC_NUM   	�INTRAC_D_T �  $INTRAC_DIV   	$�DH_EXTRA_T � 0 $VALID  $X  $Y  $Z  $W  $P  $R  �MRR_GRP_T �H �$BELT_ENABLE  $CART_ACCEL1  $CART_ACCEL2  $CIRC_RATE  $CONTAXISNUM  $PS_EXP_ENBL   $EXP_ENBL  $JOINT_RATE  $LINEAR_RATE  $PATH_ACCEL1  $PATH_ACCEL2  $PATH_ACCEL3   $PROCESS_SPD  $PROC_SPDLIM  $CNT_ACC_MGN  $DDACC_RATIO  $FWP_TIME1  $FWP_TIME2  $ACCEL_RATIO  $DECEL_RATIO  $PPABN_ENBL  $ROTSPEEDLIM  $SPEEDLIM  $SPEEDLIMJNT  $DEF_MAXACCE   $USE_CAL  $SPIN_CTRL  $SYN_ERR_LIM   $SYNC_GAIN   $SYNC_OFFSET   $MOUNT_ANGLE  $COLLINEAR  $COINCIDENT  $ACCEL_TIME1   	$ACCEL_TIME2   	$ENCSCALES   	$EXP_ACCEL   	$PS_INPOS_TI   $INPOS_TIME   	$JNTVELLIM   	$JNT23_UPLIM  $JNT23_LOWLI  $LOWERLIMS   	$LOWERLIMSDF   	$MASTER_POS   	$MIN_ACCTIME   	$MOSIGN   	$MOT_SPD_LIM   	$PERCH    	$MOVERRLIM    	$PERCHTOL    	$STOPERLIM   	$STOPTOL   	$SERVO_CTRL  $PS_SV_OFF_A   $SV_OFF_ALL  $SV_OFF_ENB   	$SV_OFF_TIME   	$UPPERLIMS   	$UPPERLIMSDF   	$TRKERRLIM  $PAYLOAD  $PS_MAX_PAYL   $MAX_PAYLOAD  $AXISINERTIA   	$AXISMOMENT   	$MAX_AMP_CUR   	$ACCEL_PARAM   $MAX_PTH_ACC  $MRRDUM2   $PS_BCKLSH_C   $BCKLSH_COUN   	$MOVER_GAIN   	$MOVER_SCALE   	$MOVER_OFFST   	$CLALM_TIME  $TSMOD_TIME  $CHKLIMTYP  $SNGLRTY_STP  $INPOS_TYPE  $JOG_TIME_M  $MIN_ACC_UMA  $MIN_ACC_UCA  $ACC_SCL_UCA  $SLMT_J1_LW   $SLMT_J1_UP   $SLMT_E1_LW   $SLMT_E1_UP   $SLMT_J1_NUM  $SLMT_E1_NUM  $PS_SPCCOUNT   $SPCCOUNTTOL   	$SPCMOVETOL   	$SHORTMO_MGN  $MIN_ACC_CMC  $EXTACCRATIO  $CN_GEAR_N1  $CN_GEAR_N2  $SFLT_ERLIM   	$SV_CTRL_TYP   	$PS_CARTMO_M   $CARTMO_MGN  $MIN_CAT_UMA  $MIN_ACC_SHM  $GEAR_RATIO   	$EXP_JOG_ACC   	$PS_ARMLOAD   $ARMLOAD   $ACC_PA_UMA  $ACC_PC_UMA  $AXIS_IM_SCL  $PS_MOT_LIM_   $MOT_LIM_STP  $JG_FLTR_SCL  $JOGACCRATIO   $TORQUE_CONS   	$MIN_PAYLOAD  $DECOUP_MGN   $DECP_MGN_WR   	$PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $FFG_MGN_J2  $FFG_MGN_J3  $DVC_AC0_MAX   	$DVC_AC1_MAX   	$DVC_ACC_MAX   	$DVC_ACC_MIN   	$DVC_JRK_MAX   	$DVC_JRK_MIN   	$SV_DBL_SMT  $SV_MCMD_DLY  $SV_GRV_X  $SV_GRV_Y  $SV_GRV_Z  $SV_DH_D   	$SV_DH_A   	$SV_DH_COSA   	$SV_DH_SINA   	$SV_LNK_M   	$SV_LNK_X   	$SV_LNK_Y   	$SV_LNK_Z   	$SV_LNK_IX   	$SV_LNK_IY   	$SV_LNK_IZ   	$SV_Z_SIGN   	$SV_DMY_LNK   	$SV_DH_COSTH   	$SV_DH_SINTH   	$SV_THET0   	$LNK23Z  $LNK23X  $LNKCBZ  $LNKCBX  $CB_MASS  $CB_IX  $CB_IY  $CB_IZ  $LNKSBY  $LNKSBX  $LNGTSB  $SPCNS  $ARMLOAD_X   $ARMLOAD_Y   $ARMLOAD_Z   $DUTY_ENB   	$DUTY_PARAM1   	$DUTY_PARAM2   	$QSTOP_TOL   	$NE_ENB  $LINK_TYPE   	$ARMLOAD_NUM   	$DH_THETA0   	$DH_THETA   	$DH_D   	$DH_A   	$DH_ALPHA   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	$DH_VD   	$DH_VA   	$DH_VALPHA   	$LINK_VM   	$LINK_VSX   	$LINK_VSY   	$LINK_VSZ   	$LINK_VIX   	$LINK_VIY   	$LINK_VIZ   	$DH_HD   	$DH_HA   	$DH_HALPHA   	$LINK_HM   	$LINK_HSX   	$LINK_HSY   	$LINK_HSZ   	$LINK_HIX   	$LINK_HIY   	$LINK_HIZ   	$DH_OTHETA   	$DH_OD   	$DH_OA   	$DH_OALPHA   	$LINK_OM   	$LINK_OSX   	$LINK_OSY   	$LINK_OSZ   	$LINK_OIX   	$LINK_OIY   	$LINK_OIZ   	$FLINK_BX   	$FLINK_BY   	$FLINK_BETA   	$SPBALANCE_K   	$SPLENGTH_0   	$SPACT_X   	$SPACT_Y   	$SPACT_Z   	$SPFULC_X   	$SPFULC_Y   	$SPFULC_Z   	$INTERACTION 1� 	$AUTO_SNGSTP  $T1T2_SNGSTP  $CART_2ND_TI  $JNT_2ND_TIM   	$LC_QSTP_ENB  $CP_CUTOFFOV  $CP_MINSEG  $MASTREV_ENB  $MASPOS_DIFF   	$INTRAC_NUM 1� 	$INTRAC_DIV 1� 	$OBS_DIST  $SV_PARAM   2$MIJNTCHKLMT  $LCHWARN_ENB  $ABC_PARAM   $MECH_MASK  $MECH_TYPE  $AXS_MAP_NUM  $AXS_MAP   	$DH_EXTRA 1� 
$AXS_COUPLE   	$PS_ROBOT_CR   $ROBOT_CRC   Q�MSK_CE_GRP_T � P $T1_USERCART  $T1_USERJNT   	$T1_CARTVEL  $T1_JNTVEL   	$T1_WARNING  �MTCOM_CFG_T �  $CNC_NO  $NORES_TIMEO  �OPWORK_T �, $SYSBUSY  $SOPBUSYMSK  $TPBUSYMSK  $UOPBUSYMSK  $INTPRUNNING  $INTPPAUSED  $INTPMASK  $OPT_OUT  $UOP_DISABLE  $OUTIMAGE   $OP_PREV_IMG   $OP_INV_MASK   $ORGOVRDVAL  $USER_OUTPUT   $PS_ENBL_ON   $ENBL_ON  $MLT_RBT_ENB  $PMC_EDT_MSK   $NOALM_MSK  $DUMMY19  \�OVRDSLCT_T � x $OVSL_ENB  $SDI_INDEX1  $SDI_INDEX2  $OFF_OFF_OVR  $OFF_ON_OVRD  $ON_OFF_OVRD  $ON_ON_OVRD  $DUMMY   H�OVRD_SETUP_T � @ $OVRD_NUM  $OVERRIDE   
$OVRD_NUM_S  $OVERRIDE_S   
 �TRACECTL_T � H $TASK_STATUS  $TRC_TOP_IDX  $TRC_BTM_IDX  $TASK_ID  $DUMMY4  �TRACEDT_T � D $EPT_INDEX  $LINE_NUM  $FILE_OFST  $EXEC_TYPE  $LINE_ST  �TRACEUP_T � @ $TRC_UPDATE  $DISP_PXNN  $DUMMY2  $DUMMY3  $DUMMY4  @�PG_CFG_T � $SUBTASKNUM  $NUM_TASKS  $JMPWAIT_UPR  $JMPWAIT_LOW  $FAST_MODE  $RCVFAIL_CNT  $WAITREL_CFG  $ACC_CTRL  $CNT_CTRL  $IGNR_PLS  $DBTB_STPTYP  $BWD_CFG  $RESUME_CFG  $IGPAUS_PRI  $MTNLN_CFG  $PAUS_RTN  $RESERVE1  $RESERVE2  ��PG_DEFSPD_T � L $AP_DEF_SPD  $AP_DEF_UNIT  $DUMMY4  $APSP_PREXE  $DLY_LASTPS    ��PING_T � 0 $TIMEOUT  $DATALEN  $NPACKETS  $DEBUG  �PIPE_CFG_T � h $ARSIZE   $FILEDATA   $SECTORS  $FORMATTER  $RECORDSIZE  $MEMTYPE  $FORMAT  $AUXWORD    ��PLID_CFG_T �  $COMP_SWITCH    D�MAX_PLD_CAL_ � $ $AA  $BB  $CC  $DD  $EE  �CALC_RESULT_ � � $PAYLOAD  $PLD_J3ARM  $INERTIA4  $INERTIA5  $INERTIA6  $MOMENT4  $MOMENT5  $MOMENT6  $COMB_LOAD4  $COMB_LOAD5  $COMB_LOAD6  $PUB_INRT4  $PUB_INRT5  $PUB_INRT6   �PLID_GRP_T �P H$PI_ENB  $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $ARMLOAD3  $ROB_TYPE  $DATA_NUM  $SPEED_HIGH  $SPEED_LOW  $DEFSPD_HIGH  $DEFSPD_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DEFACC_HIGH  $DEFACC_LOW  $SAMPLE_TIME  $SAMPLE_HIGH  $SAMPLE_LOW  $MOV_AXIS   	$MOV_POS1   	$MOV_POS2   	$MOV_DEF1   	$MOV_DEF2   	$ROT_INERTIA   	$MAX_VEL_HI   	$MIN_VEL_HI   	$MAX_ACC_HI   	$MIN_ACC_HI   	$MAX_VEL_LOW   	$MIN_VEL_LOW   	$MAX_ACC_LOW   	$MIN_ACC_LOW   	$GAMMA   	$STOP_DATA  $GETDATA_FIN  $ID_RESULT   
$CALIBRATE  $PI_DEBUG  $HIDAT_V_MAX   	$HIDAT_V_MEA   	$HIDAT_A_MAX   	$HIDAT_A_MEA   	$LWDAT_V_MAX   	$LWDAT_V_MEA   	$LWDAT_A_MAX   	$LWDAT_A_MEA   	$CALC_TYPE  $MTN_CALCTYP  $CHKER_VER $PDCK_RB_TYP  $I_FACTOR   $MAX_PAYLOAD  $MAX_INERTIA   $MAX_MOMENT   $COMB_LOAD   $MAX_PLD_CAL �$IM_SRCH_DT  $WARN_DISP  $WARN_LEVEL  $OVER_LEVEL  $CALC_RESULT �$PAMSWFLG  $AMLD_SCRN  $DUMMY69  $DUMMY70  $DUMMY71   |�PLID_SV_T �P $CUR_SCRN  $CUR_GROUP  $PS_SAVE_DON   $SAVE_DONE  $NO_RECOVER  $RESULT_SAV   
$PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $DO_DEFAULT  $MOV_POS1   	$MOV_POS2   	$SPEED_HIGH  $SPEED_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DO_DEF_POS   ��PLIM_GRP_T � � $MAX_PYLD  $AXISINERTIA   	$AXISMOMENT   	$AXIS_IM_SCL  $PS_LIM_WT_S   $LIM_WT_SCL  $LIM_INR_SCL   $LIM_MNT_SCL   $LIM_CL_SCL   $PLD_MODE  $DUMMY10  $DUMMY11   ��PLMR_GRP_T � � $PYLD_ENB  $WMR_ENB  $ANGLE  $PLMR_AA  $PLMR_BB  $PLMR_CC  $PLMR_DD  $PLST_ANG   
$COMP_SW  $MAX_XY_LOC  $MAX_Z_LOC  �PLST_GRP_T � p $COMMENT $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  �PL_RES_G_T � | $PAYLOAD  $SAVMOMENT4  $SAVMOMENT5  $SAVMOMENT6  $SAVINERTIA4  $SAVINERTIA5  $SAVINERTIA6  $EST_RESULT    ��PL_RES_V_T �  $PL_RES_G_P   �PMON_QUE_T � 8 $QCOUNT  $QTHRESHOLD  $QHYSTERESIS  $QUEUE_UP  �PM_GRP_T � � $ACC_TIME1  $ACC_TIME2  $POS_ERR_LIM  $ROT_ERR_LIM  $ENABLED  $DBG_MASK  $COMP_SWITCH  $BWD_ACC1  $BWD_ACC2  $JVEL_RATIO  $REWIND_NUM  $GTF_ACC1  $GTF_ACC2  �POCFG_T �   $PODEBUG  $OVERRUN_TOL   ��PODATA_T � P $OVERRUN_CNT  $CUR_INDEX  $PROGRAM_ID   2$LINE_NO   2$OVERRUN_ITP   2�POINFO_T �  $CUR_INDEX  $INFO   �@x�POIO_T � ( $SLEQ_NUM  $IO_TYPE  $IO_INDEX  `�POS_EDIT_T � � 	$LOCK_POSNUM  $HIDE_MENU  $HIDE_POSNUM  $AUTO_RENUM  $COPY_POSDAT  $AUTO_RENUM2  $RMV_MANRENM  $COPY_POSTYP  $CPRUT_ENB   �PRGADJ_T � h $X_LIMIT  $Y_LIMIT  $Z_LIMIT  $W_LIMIT  $P_LIMIT  $R_LIMIT  $SPEED_ADJ  $NEXT_CYCLE  \�PRGNS_CFG_T � � $ALGO_VER  $NYQ_FREQ  $WIN_TYPE  $WIN_SIZE  $OVERLAP  $FREQ_LIM  $MIN_NUM  $CREATED  $VERIFY  $PROGNAME %$CREATE_GP  $STATUS_GP  $DEBUG  $MAILTIME  $MAILEVENT  $LASTMAIL  �PRGNS_ELEM_T � � $ENABLE  $FEASIBLE  $AXIS  $PS_ELEM_NUM   $ELEM_NUM  $ROT_RATIO  $MAX_FREQ  $THRE_REL  $THRE_ABS  $DEGRAD_LVL  $DEGRAD_BASE  $DEGRAD_RATE  $UPD_DATE $BASE_DATE ׸�PRGNS_GRP_T � X $ELEM 2� $MIN_ANG   	$MAX_ANG   	$BASE_ANG   	$LAST_MOD   	$BASE_MOD   	 ��PRGNS_PREF_T � ( $GRIDLINES  $BARS_NUM  $STYLE  *�PROTOENT_T �  $P_NAME !$P_PROTO  �PROXY_CFG_T � � $LIST_PORT  $PROXY_ENB  $PROXY_SRV )$PROXY_PORT  $DIRECT_1 )$DIRECT_2 )$DIRECT_3 )$DIRECT_4 )$DIRECT_5 )$DIRECT_6 )$DIRECT_7 )$DIRECT_8 )��PF_DATA_T �   $VALUE  $GROUP  $AXIS  )��PF_CFG_T �| $ENABLE  $PROG_NAME %$CUR_GROUP  $RAN_GROUPS  $START_TYPE  $TOTAL_TIME  $TOTAL_PWR  $INS_PWR  $REGEN_PWR  $INS_REGEN  $EXE_DATE $DATA_TYPE  $RES_NAME %$MONTR_RATE  $D_PWR_SUP  $D_PWR_REG  $RV_LIM1  $RV_LIM2  $DEGREE  $REFRESH  $OVERRIDE  $RV_HRS_DAY  $RV_DAYS_YR  $MAXSIZE  $SUMMARY 2� $CONFIG_SET  $SUPPORT  $LAST_RUN  %��PF_PREF_T � 4 $GRIDLINES  $BARS_NUM  $DATA_TYPE  $STYLE  �PSSAVE_T � $MC_FOLDER 	$SLAVE_SAVE  $START_MULTI  $SLAVE_LOAD   $LOAD_DEV  $KEEP_HNADDR !$KEEP_HRADDR !$KEEP_CCOMM $KEEP_CPROT 	$PS_KEEP_COP   $KEEP_COPER  $KEEP_CSTATE  $KEEP_CREMOT $KEEP_CTIMEO  $KEEP_CSREMO $KEEP_CUNAME e$KEEP_CHPWD  $KEEP_SBMSK !��PSSAVE_GRP_T � , $FLANGE  $SYNC_FLANGE  $SYNC_MST_CN  �PS_CONFIG_T � � $DB_IMMTRIG  $DA_IMMTRIG  $DB_NOTRIG  $DA_NOTRIG  $TCLAMP_WARN  $USE_DYNSPD  $MAX_SEARCH  $NUM_PSMOTN  $DB_MARGIN  $RESOLUTION  $COMP_MASK  $PX_STARTED  $SCAN_READY  $SCAN_ALIVE  �PS_CP_CFG_T �  $ENB  $REF_MODE  �PS_CP_GRP_T � � 
$ENB  $REF_MODE  $FLANG_VALID  $FLANG_TICK  $FLANG_TRANS $PREVI_TRANS $UTOOL_VALID  $UTOOL_TRANS $FKSOL_FP  $SEG_COUNTER  L�PS_ITEM_T � � $BASE_DIST  $TUNE_MSEC  $MN_LEN  $ITEM_LINE  $ITEM_DONE  $TRIGGERED  $STOP_TRIG  $NG_ITEM  $CLAMPED  $PARAM1  $PARAM2  $PARAM3  $ML_ACT_P  $MN_CODE   �PS_MOTION_T ��  $OWNER_TID  $G0  $PS_DONE  $PG_STATUS  $DB_STATUS  $DA_STATUS  $DB_MIN_DIST  $DA_MAX_DIST  $PARENT_NAME %$CHILD_NAME %$PARENT_LINE  $SCAN_COUNT  $SEG_STARTED  $SEG_COUNTER  $SCAN_ABORT  $PARENT_EPT  $CHILD_EPT  $PRV_VALID  $PRV_DB_DIST  $PRV_DA_DIST  $PRV_VEC   $PRV_TICK  $BASE_SPEED  $DEST_VALID  $DEST_VEC   $UT_TRANS $MMR_P  $MODONE  $NEXT_MODONE  $SMH_MASK  $NUM_ITEM  $ITEM 2� 8�PWRUP_DLY_T �   $DELAY_TIME  $SY_READY   D�QSKIP_GRP_T � � $ERROR_CNT2   	$QSKP_ERRCNT   	$QSKP_CURANG  $QSKP_CURAN1  $QSKP_CURAN2  $QSKP_CURAN3  $QSKP_CURAN4  $QSKP_CURAN5  $QSKP_CURAN6  $QSKP_CURAN7  $QSKP_CURAN8  $QSKP_CURAN9  �J2RED_T � 4 $EXD_RTQ  $EXD_ITP  $EXD_PRG  $EXD_LINE  	��RDCR_GRP_T � � $RMAX_TORQUE   	$RMIN_TORQUE   	$THRES_TORQ   	$RGEAR_RATIO   	$WARN_FLG   $COMP_SW  $RESERVE   	$SPC_ITP  $NUM_EXD  $J2TH2ND  $J2RED 1� ��REFPOS11_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  X�REFPOS21_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS31_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS41_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS51_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS61_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  L�REFPOS71_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  �REFPOS81_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPSMSK_T �  $MAXREFPOSEN    �REMOTE_CFG_T � 4 $REMOTE_TYPE  $REMOTEIOTYP  $REMOTEIOIDX   ��REPOWER_T �  $FLAG  ��RESTART_T � , $FLAG  $DSB_SIGNAL  $STARTUP_CND   ��RS232_CFG_T � � $COMMENT $DEVICEUSE  $SPEED  $PARITY  $STOPBITS  $FLOWCONTROL  $TIMEOUT  $CUSTOM  $AUXTASK  $INTERFACE  $STATUS  ��RSCH_T � @ $OLD_SPEC_SW  $FREEFROMSIZ  $TARGET_DIR 	$UPDT_MAP   �RSPACE_T �� !$COMMENT $USAGE  $ENABLED  $IN_EXTERIOR  $ENTRY  $ENT_SIGN_ON  $PRIORITY  $PRIORWRK  $DOUT_TYPE  $DOUT_INDX  $DIN_TYPE  $DIN_INDX  $FRIEND_GRP  $UFRAM_NUM  $UTOOL_NUM  $MYHOLD  $LENGTH_VTEX  $FIRST_VTEX   $SECND_VTEX   $UFINV_POST $MARGIN  $WAITING  $FIRST_VTX2   $SECND_VTX2   $G2ENTRY  $G1ENT_INTR  $G2ENT_INTR  $PRE_UFRAM  $NO_USE_DI  $HOLD_REQ  $CSPACE_NUM  $CUR_TCP   $PRE_TCP   �GP_STATUS_T � @ $IN_USE  $SPACE_NUM  $PRIORITY  $STATUS1  $STATUS2  ��COM_SPACE_T �X $USE_MLT_CTN  $H_PRIORITY  $IN_CONTROL  $IN_SPACE_GP  $WT_SPACE_GP  $USE_GP  $DEADLOCK_GP  $DELAY_CNT1  $DELAY_CNT2  $GP_STATUS 2� $DOUT1_TYPE  $DOUT1_INDX  $DOUT2_TYPE  $DOUT2_INDX  $DOUT3_TYPE  $DOUT3_INDX  $DIN1_TYPE  $DIN1_INDX  $DIN2_TYPE  $DIN2_INDX  $EXT1  $EXT2  $V1   $V2   $V3   ��GP_HOLD_T � � $STATUS  $GP_MSK  $SPACE_NUM  $CSPACE_NUM  $REQ_GRP  $PS_RATE   $RATE   $INT_POS   $ACT_POS   $PRD_POS   $S1  $S2  $S3  $S4   ��RSPACEG_T � 0 $COM_SPACE 2� $GP_HOLD 2� $SPARE_INT   
t�RSPACESR_T � � $SR_ENB_TYP   $RUNNER_AXS  $HAND_LNGTH  $HAND_THICK  $FLIP_ENB  $INTFERENCE  $HAND_IF_CHK  $HANDI_TYPE  $HANDI_INDX  $SR_G1POS   $SR_G1POS_IN   $SR_G1ANG   $SR_G1ANG_JF   $SR_PRM   	�RTCFG_T � � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $RSM_RTCP  $INLINE_WRST   $TBC_PTH_CMP  $DRTCP_ENB  $LDR_SP_RATE  $LDR_RSP_RAT  $COMP_SWITCH   &$�RV_DATA_T �  $DATETIME    	$VALUE    	�RV_DATA_GRP_ �  $DATA  2� �SCR_T �	| �$ITP_TIME  $NUM_GROUP  $NUM_TOT_AXS  $NUM_DSP_AXS  $JOGLIM  $FINE_PCNT  $COND_TIME  $MAXNUMTASK  $KEPT_MIRLIM  $MAXPREMTN  $MAXPREAPL  $PRE_EXE_ENB  $NUM_SYS_MIR  $NUM_PG_MIR  $BRKHOLD_ENB  $ENC_AXIS    $ENC_TYPE    $NUM_GP_MADE  $NUM_RLIBSOC  $NUM_MOTNSOC  $DUMMY158  $SV_CODE_OPT  $SFSPD_OVRD   $COLDOVRD  $COORDOVRD  $TPENBLEOVRD  $FENCEOVRD  $JOGOVLIM  $SFJOGOVLIM  $RUNOVLIM  $SFRUNOVLIM  $MAXNUMUFRAM  $MAXNUMUTOOL  $LCHDLY_TIME  $RECOV_OVRD  $JOGWST_MODE  $JOGLIMROT  $MOTN_PC_RUN   @$RESETINVERT  $OFSTINCVAL  $FWDENBLOVRD  $TPMOTNENABL  $PREV_CTRL  $MAX_PRE_FDO  $PRE_MB_CMP  $MB_DSBL_MSK  $MB_DSB_MSK2  $SVSTAT  $UPDATE_TIME  $JG_DSBL_MSK  $NUM_PG_AMR  $MB_LD_MSK  $MOTN_LD_MSK  $MOTN_LD_MK2  $AMP_TYPE   T$CAP_AMP_DIS   T$HBK_MAP_ENB  $HBK_IO_TYPE  $HBK_IO_IDX  $PPA_MAP_ENB  $PPA_IO_TYPE  $PPA_IO_IDX  $MOTN_LD_IDX   @$DVC_DBG  $DVC_ENB  $DVC_MODE  $DVC_MODE1  $DVC_MODE2  $DVC_MODE3  $DVC_C_RATIO  $INTASK_OVRU  $DSP_TYPE  $CABINET_TYP  $NE_MODE  $PG_DSBL_MSK  $JOG_AUX_ENB  $SUBCPU  $NE_SIN_RESO  $UPDATE_MAP1  $UPDATE_MAP2  $UPDATE_FLAG   $HW_C1_TIME1  $HW_C1_TIME2  $ATR   �$UNITTYPE   �$ATRATTRIB   �$NE_CYCLE  $NECA_OVRUN  $FLTR_2_FIX  $STARTUP_CND  $DSB_SIGNAL  $LPCOND_TIME  $CHK_CH_SCTM  $F_ATR   �$F_UNITTYPE   �$F_ATRATTRIB   �$FSSB_STAT   �$CHAIN_TIME  $CHAIN_STAT  $CHAIN_RSDN  $DSP_MAP_ENB  $IDX_TBL_MSK  $PROC_CTRL  $TEMPER_LIMS   T$FSSB1   $FSSB2   $FSSBDIAGENB  $RAILACC_ENB  $SMCR_LOADED  $DUMMY159  $PS_DSP_TYPE   $DSP_TYPE2  $PRC_DSP   $PRC_CD_ID 	$MOTN_FUNC   $INTRINS_TP  $DIAG_FUNC  $TRANS_NUM   T$TRANS_MAX   T$TRANS_WARN   T$CBLCUR_MAX   T$CBLCUR_A   T$CBLCUR_B   T$CBLCUR_WARN   T$DAC_TRANS   T$DAC_CBLCUR   T$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $CE_RIA_SW  $SAFE_SPD  $SAFE_ROTSPD  $T2_LOCK_ENB  $DSB_MOINIT  $MAX_DF_LEN  $MPDT_TIMLMT  $FAST_HRDYON  $ORG_PTH_RSM  $DAC_LMT  $MULSELENB  $UPDATE_MAP3   $JCOLDOVRD  $JTPENBOVRD  $JFENCEOVRD  $FAN_ALMLVL  $FAN_WRNLVL  $HARDTYP_MAP  $COMP_SW   2$SHADOWRECS  $SHADOWTIME  $FANSTOP_TIM  $BRK_ECO_ENB  $AUTATR_STAT  $AUTO_SBRIDX  $AUTO_DSPIDX  $AUTO_ATRIDX   $AUTO_AMPINF   �$AUTO_AMPCUR   �$REGTYPE  �AX_OFS_T �  $X  $Y  $Z  ��SCR_GRP_T �� �$NUM_SEG   $NUM_PT   $ARM_TYPE  $DUMMY121  $ARM_TYPE_B  $NUM_AXES  $NUM_ROB_AXS  $NUM_RED_AXS  $WRST_AXIS_S  $WRST_AXIS_E  $SYNC_M_AXIS  $SYNC_S_AXIS  $WRIST_TYPE  $HW_STRT_AXS  $AXISORDER   	$DUMMY122  $BRK_NUMBER   	$DUMMY123  $DD_MOTOR   	$ROTARY_AXS   	$LOADRATIO   	$CONFIG_MASK  $LINK_LENGTH   $EXT_ORDER   $DUMMY124  $EXT_XYZ_MAP   $DUMMY125  $EXT_OFFSET   $EXT_LENGTH   $ROBOT_ID $ROBOT_MODEL 	$ROBOT_FILE 	$ROBOT_INT  $SV_CODE_ID $JOGLIM_JNT   	$COORD_MASK  $OP_BRK_NUM   	$DUMMY126  $USE_TBJNT  $USE_TBCART  $NUM_DUAL  $DUMMY127  $PS_TURN_AXI   $TURN_AXIS   $AXS_AMP_NUM   	$FLEXTOOLTYP  $AXS_XYZ_MAP   	$DUMMY128  $OFST 1� 	$KINEM_ENB  $DUMMY129  $PS_UPDATE_M   $UPDATE_MAP  $TORQCTRL  $DSP_NUM   	$DUMMY130  $PS_M_POS_EN   $M_POS_ENB  $M_DST_ENB  $MOVE_DST  $MCH_POS_X  $MCH_POS_Y  $MCH_POS_Z  $MCH_POS_W  $MCH_POS_P  $MCH_POS_R  $MCH_ANG   	$MCH_SPD  $DST_MIR_P  $DPOS_DST  $DST_POS_X  $DST_POS_Y  $DST_POS_Z  $DSP_ERCNT   	$PS_DEST_DAT   $DEST_DATA_P   $ROBOT_FUNC  $PROC_AXS   	$DAC_MODE  $DAC_AXMODE   	$DAC_RATE1   	$DAC_RATE2   	$DAC_RATE3   	$DAC_RATE4   	$DAC_RATE5   	$DAC_RATE6   	$DAC_RATE7   	$DAC_RATE8   	$DAC_RATE9   	$DAC_RATE10   	$DAC_LMT1   	$DAC_LMT2   	$DAC_LMT3   	$DAC_LMT4   	$DAC_LMT5   	$DAC_LMT6   	$DAC_LMT7   	$DAC_LMT8   	$DAC_LMT9   	$DAC_LMT10   	$DAC_DEBUG   $FUNC_SW   $FUNC_VAL   $ABC_ENB  $HBK_ENBL  $MV_DIAG   
$ABC_MODE1  $ABC_MODE2  $ABC_MODE3  $ABC_MODE4  $ABC_MODE5  $ABC_MODE6  $ABC_MODE7  $ABC_MODE8  $ABC_MODE9  $SAFE_JNTSPD   	$ROBOT_LABEL $DSP_NUM_FLG  $GROUP_NUM  $COMP_SW   $AMB_TEMP  $DSP_STRT_AX  $TOT_SBR_NUM  $TOT_DSP_NUM  $TOT_ATR_NUM  $TANDEM_SUB   	$DSP_ORDER   	$ATR_ORDER    $AMPINF_ORDR    $AMPCUR_ORDR    $FIX_ORNT_WR  �SERVENT_T � $ $S_NAME !$S_PORT  $S_PROTO !0�SERV_MRA_T � d $DATETIME  $ERR_CODE  $SAFETY_ST  $IMP_VEL   	$IMP_TOQ   	$ANGLES   	$DIST_TOQ   	 h�SERV_REC_GRP � p $TOTAL  $BIN_V1T1   	$BIN_V1T2   	$BIN_V2T1   	$BIN_V2T2   	$MRA_REC 1� 
$MRA_IDX  $WCA_REC 1� 
d�SERV_RV_T �  $OVER_LIMIT   	�SERV_OCCUR_T �  $ERR_CODE  $COUNTER  2p�SHELL_CFG_T � 5$JOB_BASE  $RSR_ENABLE   $NUM_RSR   $RSR1_NAME %$RSR2_NAME %$RSR3_NAME %$RSR4_NAME %$RSR5_NAME %$RSR6_NAME %$RSR7_NAME %$RSR8_NAME %$JOB_ROOT %$CONT_ONLY  $USE_ABORT  $RSR_ACKENBL  $INVERT_CHK  $UOP_SEL_STA  $RSR_ACK_PUL  $COM_TIMEOUT  $PNS_ENABLE  $SHELL_NAME %$START_MODE  $TPFWD_KAREL  $ERR_REPORT  $OPTIONS  $QUE_ENABLE  $PRODSTARTYP  $CSTOPI_ALL  $SHELL_EXT  $SEL_TYPE  $EXT_SEM1  $EXT_SEM2  $MAINT_STYL  $ISOL_ENB  $DI_CHKTRIG  $PROD_MODE  $INIT_TMO  $MANRQ_TMO  $EXTEND_ENB  $KEYSWITCH  $STARTCHKTYP  $HEARTBEATMS  $PERM_LEVEL  $TEMP_LEVEL  $USTART_FT  $START_SIG  $DO_HOME_SOP  $REFPS_PR_ID  $DIS_STRTCHK  $CUSTOM  $E_RECOV_MSK  $SET_IOCMNT  $CSTOPI_ALL2   @�SHELL_CHK_T � D $ENABLE  $RESUME  $PROMPT  $ERRPOST  $FORCE  $WARN   ��SHELL_COMM_T � @ $FUNC  $STATUS  $PARM1  $PARM2  $PARM3  $PARM4   l�SMB_HDDN_T �  $BLOB    �SNPX_ASG_T � 0 $ADDRESS  $SIZE  $VAR_NAME %$MULTIPLY  �SNPX_PARAM_T � � $TIMEOUT  $SNP_ID 	$NUM_ASG  $NUM_CIMP  $NUM_FRIF  $VERSION  $STATUS  $DISP_INFO  $MODBUS_ADR  $NUM_MODBUS  $MODBUS_PORT   P8�SSR_T � x $SINGLESTEP  $DUMMY7  $SGLSTEPTASK   &$STEPTASKNUM  $STEPSTMTTYP  $STPSEGTYPE  $BWDSTEP  $SHOWSTMTTYP  �SVDT_GRP_T �� �$DATA00   	$DATA01   	$DATA02   	$DATA03   	$DATA04   	$DATA05   	$DATA06   	$DATA07   	$DATA08   	$DATA09   	$DATA0A   	$DATA0B   	$DATA0C   	$DATA0D   	$DATA0E   	$DATA0F   	$DATA10   	$DATA11   	$DATA12   	$DATA13   	$DATA14   	$DATA15   	$DATA16   	$DATA17   	$DATA18   	$DATA19   	$DATA1A   	$DATA1B   	$DATA1C   	$DATA1D   	$DATA1E   	$DATA1F   	$DATA20   	$DATA21   	$DATA22   	$DATA23   	$DATA24   	$DATA25   	$DATA26   	$DATA27   	$DATA28   	$DATA29   	$DATA2A   	$DATA2B   	$DATA2C   	$DATA2D   	$DATA2E   	$DATA2F   	$DATA30   	$DATA31   	$DATA32   	$DATA33   	$DATA34   	$DATA35   	$DATA36   	$DATA37   	$DATA38   	$DATA39   	$DATA3A   	$DATA3B   	$DATA3C   	$DATA3D   	$DATA3E   	$DATA3F   	$DATA40   	$DATA41   	$DATA42   	$DATA43   	$DATA44   	$DATA45   	$DATA46   	$DATA47   	$DATA48   	$DATA49   	$DATA4A   	$DATA4B   	$DATA4C   	$DATA4D   	$DATA4E   	$DATA4F   	$DATA50   	$DATA51   	$DATA52   	$DATA53   	$DATA54   	$DATA55   	$DATA56   	$DATA57   	$DATA58   	$DATA59   	$DATA5A   	$DATA5B   	$DATA5C   	$DATA5D   	$DATA5E   	$DATA5F   	$DATA60   	$DATA61   	$DATA62   	$DATA63   	$DATA64   	$DATA65   	$DATA66   	$DATA67   	$DATA68   	$DATA69   	$DATA6A   	$DATA6B   	$DATA6C   	$DATA6D   	$DATA6E   	$DATA6F   	$DATA70   	$DATA71   	$DATA72   	$DATA73   	$DATA74   	$DATA75   	$DATA76   	$DATA77   	$DATA78   	$DATA79   	$DATA7A   	$DATA7B   	$DATA7C   	$DATA7D   	$DATA7E   	$DATA7F   	 8�SVPRM_UPD_T �  $PRM   
��SVGUN_CT_T � ` $OUTPUT_ENB  $INPUT_ENB  $GROUP_NUM  $AXIS_NUM  $GO_VALUE  $GI_VALUE  $IO_SCALE  �SYSLOG_T � � $SIZE  $MODE  $STATUS  $ADDRESS  $DATA_SIZE  $COMP_VALUE  $STOP_MODE  $CURR_VALUE  $FLOG_ID_LO  $FLOG_ID_HI  $FLOG_ID_IN  $FILE_OUT  $FILE_NAME $ID  x�SYSLOG_SAV_T � h $SAVE_BLCKS  $SAVE_TASKS  $SAVE_D_CPU  $SAVE_D_SIZ  $SAVE_D_ADD  $FILE_OUT  $FILE_NAME ��SYSTEM_TIMER � p 
PWR_TOT  PWR_LAP  SRV_TOT  SRV_LAP  RUN_FLG  RUN_TOT  RUN_LAP  WIT_FLG  WIT_TOT  WIT_LAP  �TBC_ACC_T �X -$ACC_LEN1  $ACC_LEN2  $ACCEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT   	$M_STAT  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $AC_ACC  $JK_ACC  $VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AAL1  $AAL2  $AAL3  $AAL4  $AAL5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM   
��TBCCFG_T � ` $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $TBC_STAT   $TC 2� $TBC_DEBUG  �TBCSG_GRP_T � \ $ENABLE  $APPRC_SCL   
$OPEN_SCL   
$CLOSE_SCL   
$CLS_MINF2   
$CLS_MINACC   
�$$CLASS  ������       �$$VERSION  ������  ���$AAVM_WRK 2 ������ 0  �5�                                �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            XMOD�                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            $OR�                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            DYN_�                                                 	 	                                     ���� 	                                     ����                                                       	                                                             �$ABSPOS_GRP 1������� <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �$ACC_MAXLMT         ��   ��$ACC_MINLMT        ��    �$ACC_PRE_EXE        ��    �$AC_UPDATE  �����������$ALARMRECOV ������   �        �$ALMDG ������                �$ALM_IF ������    d                                                                                                       d                                                                                                         , 
                                         �$ANGTOL  ������� 	 A   A   A   A   A   A   A   A   A   �$APPLICATION ?������� 
 HandlingTool          
V8.20P/A2          x.p
88150              80 
3348966            xis
91                 pra
V8.20P/A2          rod7DE3/A2            pc 	80604.015          Y pFRL                ld32                  V��$AP_ACTIVE      ����   �$AP_AUTOMODE         �    �$AP_CHGAPONL         �   �$AP_COUPLED 1�������                                                                  �$AP_CUREQ 1������   T                                          	           	            	 ���                                          	           	            	 ���       �Handling      HT           	           	HTTHKY     	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ����$AP_CURTOOL      ����   �$AP_DO_CLEAN         �    �$AP_DO_CLENM  �������                                                                                                                          �$AP_DSPDRYRN         �    �$AP_HIDE  ������� @                                                                                                                                                                                                                                                                 �$AP_MAXAPP         �   �$AP_MAXAX          �    �$AP_PLUGGED      ����   �$AP_PRC_DSBM  �������                                  �$AP_PROC_DSB         �    �$AP_SEGF_CHK         �    �$AP_SEG_CHKM  �������                                                                                                                          �$AP_SELAP  ������� @                                                                                                                                                                                                                                                                �$AP_TOTALAX      ����    �$AP_USENUM  �������   �$ARG_STRING 1������� 
�MENUS             
MENU_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                I/O SIGNALS       Tryout Mode       Input Simulated   Output Simulated  OVERRIDE = 100    In cycle          Prog Aborted      Tryout Status     	Heartbeat         MH Fault          MH Alert            n                  n                  n                  n                  n                  n                  n                  n                  n                  n                TOOL              
TOOL_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                WORK              
WORK_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                POS               	POS_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                DEV               	DEV_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PALT              
PALT_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                GRIP              
GRIP_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                USER              
USER_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PREG              
PREG_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                �$ARG_WORD ?	�������  	$         	[         	]         	�          	�          �$ASBN_CONFIG �������           �$ASCII_SAVE            �    �$ATCELLSETUP 	�������%  OME_IO                               %MOV_HOME                              %MOV_REPR                                      �$AUTOBACKUP 
�������    FRA:\                                             '`                       �                 15/12/03 07:34:46         �                          �                          �                          �                            ��                                                                                                                                       ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      �  RA:\_BACKUP_\ATBCKCTL.TMP DATE.DT                                                                                                �$AUTOINIT         �    �$AUTOMESSAGE        �   �$AUTOMODE_DO         �    �$AUTOMODE_OV         �   �$AUTOPAUSPOS !��������  (7����������������������������)����������������������������9����������������������������I����������������������������(O����������������������������(O����������������������������(O����������������������������(O�����������������������������$AUTOPPOSTSK  �������                                  �$AUTOUPDTMOD         d�   �$AXIS_COUNT 1������   �  � 	  �@�_�Aw �� �^� *58             	  VJ z�` Uj `�  Z�o ?�~             	                                      	  U�p ��H���j�����V�             	                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXIS_METER 1������   �  P 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXSCRDCFG 1������  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �$BACKGROUND         �   �$BACKUP_NAME 	�������	BACKUP    �$BACK_EDIT 1������� 
 �%-BCKEDT-                              %FOLGE011                              �     ��%-BACKUP-                              �    �                        %-BCKEDT-                              ��%-BCKED2-                              %                                       	L       %-BACKU2-                                    �                        %  BCKED2-                              ��%-BCKED3-                              %UP001                                        %-BACKU3-                                    �                        %-BCKED3-                              ��%-BCKED4-                              %                                       	��      %-BACKU4-                                    �                        %-BCKED4-                              ��%-BCKED5-                              %�                                      ���      %-BACKU5-                                    �                        %-BCKED5-                              ��%-BCKED6-                              %�                                      ���      %-BACKU6-                                    �                        %-BCKED6-                              ��%-BCKED7-                              %�                                      ���      %-BACKU7-                                    �                        %-BCKED7-                              ��%-BCKED8-                              %                                       ���      %-BACKU8-                                    �                        %-BCKED8-                              ��%-BCKED9-                              %                                       ���      %-BACKU9-                                    �                        %-BCKED9-                              ��%-BCKCRT-                              %�                                      ���      %-BACCRT-                                    �                        %-BCKCRT-                              ���$BCK_NO_DEL         �   �$BGE_UNUSEND         �   �$BLAL_OUT �������  �   �$BWD_ABORT         �    �$BWD_ITR_RTN         ��   �$BWD_NONSTOP         �   �$CE_OPTION         �   �$CE_RIA_ID         �   �$CFCFG �������                      �$CF_PARAMGP 1�������                                                                                                     C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  C�  D  D  D  D  D    C�  C�  C�  C�  C�  C�  D	� D  D"� D/  D;� DH  DT� Da  Dm� Dz  D�@ D�� D�� D�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�  �$CHECKCONFIG         �    �$CHG_PRI 1�������         ��������������������������������������������������������������������������������������������������������������������$CHKPAUSPOS 1�������  ,    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    �������������������������������$COCFG �������              �$CO_MORGRP 2�������  �   B�)�?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  �$CO_PARAMGRP 2�������  ,       ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�  �$CPCFG ������          a�-                                                                                   
                                            ����                @                                 �`        �$CPDBG ������        )cpmidbg                                      �   �  :�  7}  7~       )cpmpdbg                                      �     �  	u  	v       )midbg                                        �     �  d  e       )mpdbg                                        �     �  e  f       )mgdbg                                        �     �   Y   Z       )mfdbg                                     ���������                    )ud1:                                              �$CPDBGDEF ������       )ud1:cpdbgbuf.txt                             �                    �$CP_L64FIX ������                                                                                                                                                                                                                                                                                                                                                                                                                                               �$CP_MCRGRP 2������     d   d   d   d   d   d   d   d   d   d   d   d�$CP_MORGRP 2������  �                 >�5�CH  BH   	 B��/B���B��`B�TGB�ԩC12�             	 D*��D:hAC�0�D��DL�QDi]h             	 E���F.I�E�wF.��F&"�F:�            ?�                              CH  BH   	 F �S                                 	 IQ7                                 	 M5'                                ?�                              CH  BH   	 F�W                                 	 IJ�T                                 	 M�$                                ?�                              CH  BH   	                                      	                                      	                                     ?�         �$CP_PARAMGRP 2 ������ <                        �  �     �  x    	 C>  C>  C>  C�  Cp  D>               	 D>  D  D��fE�  D�  Em�              	 D�  Dz  EC  F�  E��fE��f            ?�  >�33 ;��?   ?�         n   @   @�   5�@333@   ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    �������$CP_RSMOFST ������                  �$CP_T1_MODE !������     G   
?@      ;��
                                               �$CP_TESTDEF ������           �$CRCFG "�������                             C4  A�             �   x   A�  Cz  B�  CH  B�  CH  C  @�     -       :d�
�$CRI_CFG #�������   �$CRT_DEFPROG %�������%�                                      �$CRT_INUSER         �    �$CRT_KEY_TBL  ������   	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������͓�����������������������������耇���������������������$CRT_LCKUSER         �    �$CRT_USESTAT         �    �$CR_AUTO_DO        ��    �$CR_INDT_ENB         �   �$CR_T1_DO        ��    �$CR_T2_DO        ��    �$CSTOP         �   �$CSXC_PARAM 2$������ 
 8
SONY XC-56                    �  �@���?�     ( АSONY XC-HR50                  �  �@���?�     ( АSONY XC-HR57                  �  �Aff?�     ( А�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �$CTRL_DELETE         �   �$CT_POPUP             �    �$CT_QUICKMEN         �    �$CT_SCREEN �������kcsc  �$CT_USERSCRN �������c_sc  �$CUSTOMMENU 1%������  <               %                                                          %                                       ���               %                                       ����              %�                                      ����              %�                                      ���Start SM Comm %IBSCMANS                              ���End SM Comm   %IBSCMANE                              ���User Cancel   %UCANCACT                              ���
User Reset    %URESACT                               ����              %�                                      ����              %�                                      ����              %�                                      ���Zange         %ZG_MENUE                              ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���VAG_KONFIG.   %VW_MENUE                              ����              %�                                      ���VAG-Dateien   %DATEIEN                               ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���
Macro Step tt %MSK_STAT                              ���Wait Monitor  %SHTPEST                               ����              %�                                      ����              %�                                      ���CYCLE POWER   %PWDCYCLE                              ���
POWER DOWN    %	PWD_MAINT                             ����$CUST_MANUAL         �   �$CZCDCFG &�������            	                                              ?|(��$DBCONDTRIG         �   �$DBLOVRD_ENB         �   �$DBNUMLIM        d�   
�$DBPXWORK 1'�������                                                                                                                          �$DBTB_CTRL (�������                ���$DB_AWAYTRIG      GCP �=��
�$DB_AWAY_ALM         �    �$DB_CONDTYP         �   �$DB_DBG 1)�������  , 
               	�       	X  	W        
                                        �$DB_MINDIST      GCP �@�  �$DB_MONTIME        ��  ��$DB_MONTYP         
�   �$DB_MOTNEND         �   �$DB_RECORD 1/�������  �                        G�O�G�O�   #            U�UY    U�EXECUTING

 ��2                                                                  G�O�                                    G�O�G�O�   $            U�UO    U�EXECUTING

 W0�                                                                  G�O�                                    G�O�G�O�               U�UI    U�EXECUTING

 �d �                                                                  G�O�                                    G�O�G�O�               UU�          XECUTING

 0 b#                                                                  G�O�                                    G�O�G�O�   	            UcU
          CANCELLED
 �0�                                                                  G�O�                                    G�O�G�O�               U�U�    U!EXECUTING

 �/��                                                                  G�O�                                    G�O�G�O�                                  XECUTING
������                                                                  G�O�                                    G�O�G�O�                                  XECUTING
������                                                                  G�O�                                    G�O�G�O�                                                ���                                                                G�O�                                    G�O�G�O�                                                ���                                                                G�O�                                    G�O�G�O�                                                ���                                                                G�O�                                    G�O�G�O�                                                ���                                                                G�O�                                    G�O�G�O�                                                                                                                   G�O�            �$DB_TOLERENC      B�  �=L���$DCSS_DEVICE 10������                                                                                                                                                                                                                            �$DCSS_LS 11������                                                                                                                                                                  �$DCSS_PARAM 2������                 �$DCSS_RBT 24������ 8 
 <                  Cπ       �   �H       �H                       Cg        ��  ��  �\  �g@ ��  �\                    C��       ��  B   ´                                B�                �z          ă@                   C1            �  B�      �  ��         c                                                     c                                                     c                                                     c                                                     c                                              C�y�Dz  C�9�Dz   	 A���A�ffAI��A;33Ad  A�               	 B�  B�  B�  B�  B�  C>               	 BffB��BffB-��B*ffB�               	 B�  B�  B�  B�  B�  C>               	  }<� �b� K�@ P   P   P                   
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                         �$DCS_CFG 5�������          dMC:\DCSL%04d.CSV                     c                   �    A   A   CH  Cz                                                                                �            �   �   �   �   �   �   �            �`iMU��    �$DCS_CRC_OUT 6�������                  �$DCS_C_FSI ?������ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_FSO ?������ P �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_RPI ?������  �                      �                      �                      �                      �$DCS_C_RPO ?������  �                      �                      �                      �                      �$DCS_SGN 7�������,�0�12-JUN-24 17:05   ���03-DEZ-15 07:35            IX�SIX�SH-�H-�                    ,�0�G���i�ZX�_                  �$DCS_VERSION �������V3.3.2            �$DEFLOGIC 18�������  	�          ���	�          ����	�          �����$DEFPROG_ENB         �   �$DEFPULSE         ��   �$DEF_ACCLIM        ��   ��$DEF_WRSTJNT         �����$DEMO_ENB            �    �$DEMO_INIT 9���������������� ���$DEMO_OPT_SL ?	������   � 
 	R575      	R745      	R746      	R747      	R750      	R751      	R752      	�          	�          	�          �$DEMO_OPT_TO  ������   � 
                                         �$DEV_INDEX         d�   �$DEV_PATH A�������A\KJLTVL111180R01\ 01\  \ \ 80\  H\ UN\ H\                         �$DHCP_CLNTID ?�������  �                  �                  �$DIAG_GRP 2>������ �    	 E�  F,D F,D E(p E(p D�               	 B�  B�  B�  B�  B�  B�               	 B�  B�  B�  B�  B�  B�               	 CeEC�  C��CG�SCEZXB�Gm            f362 678901234567890          �  A���A�=qA�A�33A�z�A��A��RA���A�=qA���                  @�  A   Ap  A�  A�  A�  B  B   B4                        ������       
  A�A�{A�=qA�=qA�{A�A�G�Aď\A��A�Q����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A�=qAυAʣ�AŮA��\A�G�A��A�ffA���A��R���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A_�AZffAUG�AO�
AJ=qAD��A>�RA8��A2ffA,  ���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A`��A[�AV{AP��AK
=AE�A?33A8��A2�\A+�
���������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A��
A��RA
=Axz�AqAj�RAc�A\Q�AT��AL�����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
 	 A�z�A�{A��\AJ=qAK
=Aq             	 =�G�=�G�=�G�>8Q�>8Q�>8Q�             	 8��b8��b8��b7�Ŭ7�Ŭ7�Ŭ             	 @ʏ\@ʏ\@ʏ\@�p�@�p�@�p�              @�  Ah  A�       	 <�C�<�t�=�P=�hs=�t�=��P             	 ;��
;��
;��
<#�
<#�
<#�
                 �?+ƨC�  <(�U     4 	 @���@���@���@���@���@���            A@     ?     	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	 ?Tz�?Tz�?Tz�?#�
?#�
?#�
             	 ��G���G���G���G���G���G�             	 B   B   B   B   B   B                	 Bx  Bx  Bx  A�  A�  A�               	 Ce
C�  C�
CG�{CEY�B�G�             	                                	   p  �  �  p  p  p             	 Ap  Ap  Ap  Ap  Ap  Ap               	 ED  E�� E�� D�� D�� DD               	                                         8����?|uB��#?N�s>)�x?��?PP;�,ƿR�C���D	��D���   0        	                                      	                                      	                                  C���D	��D���Cv�@�_�B�.�     	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                 �$DICT_CONFIG ?�������          eg      ���$DISTBF_TTS         
�   �$DISTBF_VER        
�   �$DMAURST         �    �$DMSW_CFG @������               �$DOCVIEWER A������     	 ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  �$DPM_CFG B������                          
        �$DPM_SCH 2H������ 
�   Schedule 1            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 2            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 3            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 4            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 5            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 6            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 7            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 8            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 9            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 10           �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz  �$DPM_SIM 2I������                                                                                                                                                          �$DRC_CFG J�������!�                                  !�                                  !�                                  !�                                  !�                                     �$DSBL_FAULT K�������        �$DSBL_GPMSK         ��    �$DTDIAG L������            UD1: 678901234567890                         P                                                                                                                                                                                                                                                                                                                                              �               @   �$DTRECP L������            
UD1:                                          P                                                                                                                                                                                                                                                                                                                                              �               @   �$DUMP_OPTION  �������    �$DUTR_CFG      ����   �$DUTR_CPMES      ����   �$DUTY_TEMP  È�3B�  �A�  �$DUTY_UNIT         �    �$DYN_BRK M�������        �$ED_SIZE    '   �  x �$ED_STATE         �    �$EMGDI_STAT      ���     �$ENC_STAT 1N������  �                                                                     
                 d                                                                                                                                                                                                                                                                                                                                                                                                                                 ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        �$ENETMODE 1O�������                                            �$ERROR_PROG %�������%�                                      �$ERROR_TABLE  �������  �������������������������������������������������������������$ERRSEV_NUM       ��   �$ER_AUTO_ENB         �    �$ER_NOAUTO P�������          *�  *�  *�  *�  *�  +                                                        �$ER_NOHIS         �    �$ER_NO_ALM 1Q�������  �         *�  *�  *�  *�  +                                                                                                                                            �$ER_OUT_PUT 2R�������    @�                ����$ER_SEV_NOAU  �������                 �$ETCP_VER !�������!�                                  �$EXTLOG_REQ        ��    �$EXTLOG_SIZ        ��    �$EXTSTKSIZ        ��  ��$EXTTOL      Dz  �A   �$EXT_BWD_SEL         �    �$EXT_DI_BWD S�������                  �$EXT_DI_STEP S�������                  �$E_STOP_DO        ��    �$FACTORY_TUN         d�    �$FDR_GRP 1T������  d 	                             	 �[���N8�T&hB�( ��� ��� ��� 	                                      	 C�_CC#1C��C�dB��B��             	 A�
Bs�B�A���A�AQ�\             	 A�(                                 	                                      	 A��A�eQB�A�v�A���Am9�             	 ���7��O������ S�
���v             	 <`�><`�><`�>                         
 FA�Bs�<`�>    B��                                          	 E�  F,D F,D E(p E(p D�               	 ED  E�� E�� D�� D�� DD               	 C��NC��NC��NB�ƈB�ƈB�ƈ             	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	 E�� E�@ E�@ E�� E�� E��              	 OHcGPPL�uSL�uSK�y
             	 ?�  ?�  ?�  ?�  ?�  ?�               	 :G:�:G:�:G:�9{��9{��9{��             	 ��s P� ��:����#��%�*             	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FEATURE U������   HandlingTool          allyEnglish Dictionary    , PaMulti Language (GRMN) t\ir4D Standard           prodAnalog I/O            VLOAAngle Shift           l.pcAuto Software Update  \pk4Automatic Backup      irpkBackground Editing    roduCamera I/F            LOADCnrRndImp             .pcCommon calib UIF      pk4dCondition Monitor     rpk4Control Reliable      ductData Acquisition      AD pDiagnostic log        
PCVDocument Viewer       wc.pDual Check Safety UIF D prEnhanced User Frame   ENDIExt. DIO Config       NDIFExtended Error Log    pk4dExtended User Frames  ckToExternal DI BWD       INT FCTN Menu Save        l, PFTP Interface         ct\jGroup Mask Exchange   VLOAHTTP Proxy Svr        pr.pHigh-Speed Skip       pkcsHost Communications   uct\Hour Meter            OAD I/O Interconnect 2    .pcIncr Instruction      csgeKAREL Cmd. Language   ct\jKAREL Run-Time Env    AD pKernel + Basic S/W    
PCLicense Checker       etwpLogBook(System)          MACROs, Skip/Offset   .pcMH Core               prngMechStop Protection   rosiMirror Shift          p.fdMixed logic           ted Mode Switch           93 RMotion Diag. Core     R808Motion Optm. Core     ng JMotion Profiler       t IIMotion logger         0\tpMulti-Tasking         prodPCM function          IF OPosition Registers    
IFPrint Function        ELSEProg Num Selection    oadiProgram Adjust         ParProgram Shift         \j76Program Status        OAD Program Viewer        DIF RDM Robot Discovery   imarRemote Conn Standard  ! prRobot Servo Code      !
ISNPX basic            596 Shift Library          H55Shift and Mirror Lib  RINTSocket Messaging      xy STCP Auto Set          prodTCP/IP Interface      1
PTMILIB Interface      .vrTP Firmware           j755TP Menu Accounting    
!
TPTX                  R558Telnet Interface      55 (Tool Offset           II) Torque Simulator I/F  tphcTouch Panel           oducTrouble Diag. & Prev.  j75USB port on iPendant  P
!Unexcepted motn Check 9 R8User Frame             "LoVCalibration Common   I) "Vision Core           phcdVision Library        ductVision SP CSUI        dhcpVision SP CSXC        EMAIWeb Plus              DER Web Server            
PRWeb Svr Enhancements   EnhiPendant              CVLOiPendant Grid Display tioniPendant Setup        d
!iRCalib. Standard     
!
iRCalibration AAVM    R558Independent Axes      77 (Independent Axes      TXPLIndependent Axes      HCSBR-2000iB/210F         b\hcAscii Program Loader  !
!Ascii Upload          d
!AutoMode TP operation 0 H5Basic Remote TCP      551 CE Mark               g R7CPRUT                 ) "CRT/Keyboard Manager  \tptCntrl stop by E-Stop  roduCollision Guard       CVLOCollision Guard Pack  ib.pConstant Path         td\tCornerDistance        .fdCycle Time Priority   ent DCS Joint Speed check  H54DCS Safe I/O connect  49 RDHCP                  
PRIDomain Name Serv.     775Dyn Path Modifier     10iAEnhanced Dry Run      D prError Code Output     1
TExt Path Optimization tm "Extended Axis Control fd
External mode select  MS
FRL Params            "LoaHMI Device (SNPX)     PartIntegrated PMC        h772Internet Conn/Custo    proJnt Position output   #1
KAREL                 773.Multi-Group Motion    ORDEOperation logbook     773 PC Interface          
TXPROFINET I/O          "AM0PROFINET Safety       773\PROGRAM/JOG Override   ! hPassword Protection   R MaPathSwitch             H80SNTP Client           LR MTCP SPEED OUTPUT      
TXUser Function         "LRHUser Socket Msg       801\VAG Package            ! hVAG servogun setup    R MaVAG setup 3            H80Weaving               LR MiRCalibration VAxis   
TX64MB DRAM             "LR564MB FROM             802\Arc Advisor            ! hAux Servo Code        R MaCell I/O              09
Common shell          MateCommon shell core     OAD Common softpanel       #1Common style select   lr2cCorner Region         9.fdCycle time Opt.        200DCS Pos./speed common 
PRIDisp 2nd analog port  e 20EMAIL Enhancements    OAD Email Client           #1Enhanced Rob Serv Req lr5aEnhanced T1 Mode      8.fdExt weave sch          200Extended Axis Speed   
PRIFunc stup             e 20OPT TP Ins            OAD PC Send Macros         #1Real Simple Syn.(RSS) lr5lRequires CP           0.fdRobot Library Setup   ate Robot Service Request 
PRISMB Client            MateSSPC error text       OAD Soft Limit             #1Space Check           h681TCP Speed Prediction  L
!TCPP Extention        LoadTrack Instruction     iA/5Tracking Softpart     roduVAG Software          ENDIistdpnl               fd -VAG V8.x Customizatio DER VAG EMZ & EQ Tools    5 (LFREU late Updates     
TXUpdate VAG PMC        "LR2Ascii Upload when arg 755\Profinet and CD Setti D pr*.pc protection and u ENDIDryR.Skip PWF,VAGBCK  fd -Activate CD Setting   d MoVAG Menu to Page 1    686 Implement Feedb.Tig/T 9 (CFix upper limit of GO II) To fix skip problem   sfmnFiles Updated         oducActivate CD-PS-Impr   LOADDiff.a.DryS.PN:FW-CHK JG" Diff.a.DryS.PN:FW-CHK \cdcCD:Fix SSTEP and BWD  roduFix.Er.after 8xVag_C. ! j6Update several Issues ick Enh.Alloc.Mem.CD-Mot  629To fix skip problem I ick Fix Err.Karel Var.Scr XPLOFix DCS FB_CMP alarm  MNSTFix overwr.VAG FUNC-M !
!Restore Optimizations RDERFix.Karel User n.save 65 (ZIP cmd.er.handl.impr D prRestore Optimization   #1VAG Sign Off Function funcATSHELL Heartbeat Opt 
!
No Outp.On/Off w.SRVO  ProFix-PS strt move away 6 H5GunM.DO.Prot.Gen.Opt. R716Fix iPend.scrn freeze art P381+Investig.Patch   eldpFix ABC Over Run      VLOAOver.disp.unexp.clear gex.Inv.probl.about PGPX  procRes.TCPspdoutVar E-St oducFix ABC Ov.load MSTP  PCVLModification of iRCal 3wp0Unzip Inst+Improv.    ldprFix PGPX OX-144 probl prodEnh.DryRunP.Canc/Res  
PCFix OS144 Motn-UserCa psg.Improve VAG-Backup    
!Improve VAG-Backup     Anl�                      R788�                      rc W�                      ) "�                      anlg�                      uct\�                      AD p�                      IF  �                      fd -�                      
IF �                      8 J6�                      (Lin�                      I) "�                      o\aw�                      prod�                      PCVL�                      ealk�                      leco�                      wmle�                      MH C�                      48 H�                       MHC�                      TXPL�                      d "F�                      \mht�                      PLOA�                      "APF�                      htoo�                      OAD �                      ETU"�                      ool\�                      \mht�                      tool�                      ol E�                        ��                      fdcs�                      uct\�                      PCVL�                      r
E�                      545.�                      
IF�                      73 H�                      H574�                      45 (�                      I) "�                      pfat�                      duct�                      j545�                      cens�                      CHK �                       H54�                      RINT�                      Chec�                       pro�                      VLOA�                      r
E�                      h550�                      ORDE�                      96 H�                      H552�                      50 (�                      TXPL�                      "MNA�                      550\�                      D pr�                      F  !�                       Mul�                      J600�                      6 H5�                      552 �                      0 (M�                      
TX�                      l "M�                      d
!�                      ic
�                      90 H�                      H551�                      ng J�                      I) "�                      sfmn�                      oduc�                      
EN�                      tlog�                      
!�                       H57�                      51 H�                       R54�                      art �                      xtlo�                       ! e�                       - V�                      ER V�                      H558�                      2 J8�                      (Vis�                      
TXP�                      is "�                      l.fd�                      lib.�                      RCL �                       H54�                      52
�                      alib�                      TXPL�                      vm "�                      t\cv�                      TXPL�                      ft "�                       Tt�                      igna�                      D pr�                      " #1�                      etac�                      oduc�                      CVLO�                      ta.p�                      \cb_�                      t\cb�                      rodu�                      
PC�                      lear�                      cbsi�                      rodu�                      
PCV�                      adsi�                      sig\�                      rodu�                      VLOA�                      rr.p�                      \cb_�                      t\cb�                      rodu�                      
PC�                      unsi�                      sig\�                      rodu�                      CVLO�                      ftn.�                      g\cb�                      duct�                       cbs�                      a Ac�                      631 �                       H55�                      CO R�                      RRS2�                      4 FC�                      009 �                       R58�                      631 �                      II) �                      tdme�                      duct�                      rodu�                       pro�                      AD p�                      IF  �                       MAC�                      ORDE�                      51 H�                      SEND�                      3 RR�                      551 �                       J98�                      MACR�                      ) "�                      mnmc�                      uct\�                      XPLO�                      ACR"�                      3\sf�                       H56�                      \j50�                      F
T�                      of "�                      t\j5�                      ORDE�                      oduc�                      NDIF�                      ol.f�                      ER H�                       (Fl�                      �)��                      iB/2�                       pro�                      
TX�                      t "H�                      d
!�                      10F�                       "Lo�                      F, P�                      ct\h�                      OAD �                      1" #�                      strb�                      \h60�                      rodu�                      LOAD�                      c
I�                      oduc�                      
END�                      arm.�                      RDER�                      50 (�                      IF O�                       R65�                      G.$P�                      
EN�                      frlp�                      IF O�                      g R6�                       "
�                      RDER�                      YSCF�                      NDIF�                      
EN�                      j507�                      
IF �                      3 H5�                      574 �                      7 (P�                      "
T�                      t "T�                      \j50�                      F  !�                       Inc�                      ER J�                      H558�                      1 H5�                      J510�                       II)�                      \sfm�                      j510�                       Met�                      1 H5�                      548 �                      oadi�                      t II�                      3\mn�                      prod�                       ! j�                      osit�                      ER J�                      H596�                      8 H5�                      ding�                      s, P�                      ct\j�                      PLOA�                      NPR"�                      
! �                      
!�                       H57�                      51 H�                       J51�                      II) �                      ���                      prod�                      1
T�                      cf "�                      t\j8�                      rodu�                      LOAD�                      
PC�                      nit.�                      \plc�                      !
!�                      ion �                      1
P�                      e Ge�                      
TXP�                       "K2�                      r674�                      AD p�                      " #1�                      ngcr�                      duct�                      PCVL�                      t.pc�                      ngda�                      674\�                      duct�                      AD p�                      
PCV�                      i2.p�                      sngc�                      674\�                      ct\r�                      rodu  H552  ec.pH521  AD pH532  674\R782  c
PH550  roduJ614  sngpATUP  CVLOJ545  ct\rJ616  us.pVCAM  AD pCRIM  674\CUIF  
PCVJ628  ductCNRE  at.vR631    ! RSCH  
!
DOCV  d - DCSU  ip
J604  DER EIOC  INT R542   J92R696   SkiESET  II) J516  AD pJ716  921\MASK  K207PRXY  PLOAJ627  t\j9HOCO  s "TJ513  
PCVJ542  ductJ510  skmaJ650  CVLOJ539  ct\jH510  kcklLCHK  LOADOPLG  \j92J503  r
EMHCR  j921MCSP  ! j9J506  KAREJ554  rt FMDSW  IF OMDCO  1
POPCO  adinMPRO  KARER637  rt FJ600  t IIPCMF  LOADJ514  \j97J507   "K2J515  TXPLJ517  uct\J505  209 PRST  1
TJ697  roduFRDM  kckrRMCN  " #1H930  D prSNBA  71\kSHLB  TME"SMLB  LOADR636  \j97J520  in.pHTCP  AD pTMIL  971\R789  pc
TPAC  prodTPTX  \krcTELN  
PCJ509  oducJ882  rcfcR781  PCVLJ958  uct\J957  f.vrUECK  D prUFRM  71\cVCCM  ENDIVCOR  1.fdVIPL  735.CSUI  EL UCSXC  UIFWEBP  RDERHTTP  RINTR626  g J7CGTP  L UsIGUI  IF, IPGS   "
IRCL  prodJ888  \atkH895  8" #H895  AD pH895  735\H601  K209R796  PLOAR507  t\j7J698  �9�R657   "COJ618  IF OJ858  0 H5J535  OAD J570  j670R534  "FSGJ684  NDIFR663  ER HR748  
TXJ523  oducJ555  ftpsJ568   #1R526  TXPLJ755  uct\R739  tun J985  1
TJ527  roduJ829  sgtpJ518  " #1J569  D prR651  70\sR553  979"J760  ORDER558  573J966   proR632  0\sgJ601  AT" J695  F
IR641  H590J930  XPLOJ931  ct\jJ579  57 "J541  
ENJ693  LOADR610  \j67J694  b.pcJ986  D prR648  70\sJ658  c
PJ653  roduJ656  tdflJ504  
PCVJ996  ductD064  smchF064  CVLOR666  ct\jSVMO  men.CLIO  OAD R645  j670CMSC  p.pcCMSP  D prSTYL  70\sR654  c
PCTOP  roduDCSC  sgmvR528  
PCVJNN8  ductJNN7  mkunORSR  CVLOR680  ct\jJ881  lwtpEXTS  LOADFCSP  \j67OPIS  tp.pSEND  AD pR679  670\CPRQ  .pcRLCM   proSRSR  0\swR677  c
PETSS  roduSLMT  svglJ609  PCVLJ524  uct\TCPE  iaseTOAW   ORDTRAK  H573FVAG  D prIPNL  70\sVAG1  pc
EZEQ  F ORUPD3   H57PMC3  AD pP137  670\E001  .pcE002  IF OE003  0 H5E004  OAD E005  j670E006  2.pcP170  
IF P171  90 HE007  LOADRT22  \j67E008  al.pE009  
IFP208  590 E010  VLOAE011  t\j6RT23  tol.P213  F
IP225  H590P230  CVLOP231  ct\jE013  ksevP238  IF
P244   H59E014  PCVLP246  uct\S300  kkskP275  DIFP276  R H5E015  
PCVP381  ductP477  hkkrP501  NDIFP525  ER HP537  
PCP333  oducE016  gkdfP307  ENDIP576  DER P604  3
PE018  roduP623  sgktF001  
ENDF002  RDER�      73
�      prod�      \sgk�      
EN�      ORDE�      573�       pro�      0\sg�      c
E�       ORD�      H573�      D pr�      70\s�      pc
�      F OR�       H57�      AD p�      670\�      .pc�      IF O�      0 H5�      OAD �      j670�      g.pc�      
IF �      90 H�      LOAD�      \j67�      tl.p�      
IF�      590 �      VLOA�      t\j6�      hst.�      F
I�      H590�      CVLO�      ct\j�      ftsk�      IF
�       H59�      PCVL�      uct\�      n.vr�       4$�         �      XPLO�      ct\c�      ak95�       #1�       pro�      orcm�      "CCF�      CVLO�      ct\c�      accd�      PCVL�      uct\�      pacc�      
PCV�      duct�      \pac�      
PC�      oduc�      m\pa�      c
P�      rodu�      cm\p�      pc
�      prod�      rcm\�      pc
�      prod�      rcm\�      .pc�       pro�      orcm�      t.pc�      D pr�      lorc�      sk.p�      AD p�      olor�      tsk.�      OAD �      colo�      runc�      LOAD�      \col�      csub�      VLOA�      t\co�      ccce�      CVLO�      ct\c�      acct�      PCVL�      uct\�      pacc�      
PCV�      duct�      \pav�      
PC�      oduc�      m\pa�      r
P�      rodu�      cm\p�      vr
�      prod�      rcm\�      
END�      lorc�      
! p�       - P�       Dia�      
!�      R R5�      T "L�      589 �      ol D�      cs, �       "
�      prod�      ag\p�      925"�      LOAD�      \pad�      26 "�      
TX�      oduc�      \pad�      E" #�      AD p�      adia�       "DG�      PCVL�      uct\�      adgs�      PCVL�      uct\�      mons�      PCVL�      uct\�      adgr�      PCVL�      uct\�      avrp�      PCVL�      uct\�      gse.�      OAD �      padi�      vr
�       pad�      !
!�      fd -�      e Di�      s
!�      ER R�      NT "�      R823�      se D�      cs, �       "
�      prod�      ag\s�      925"�      LOAD�      \sld�      26 "�      
TX�      oduc�      \sls�      G" #�      AD p�      ldia�       "ST�      PCVL�      uct\�      ldgs�      PCVL�      uct\�      mons�      PCVL�      uct\�      ldgr�      PCVL�      uct\�      lvrp�      PCVL�      uct\�      ldtf�      PCVL�      uct\�      edg.�      OAD �      sldi�      vr
�       sld�      !
!�       - P�      djus�       ORD�      H541�      73 H�       H54�      551 �      2
P�      adin�      Prog�      st, �       "
�      prod�      \atk�      0" #�        ��      ���      
IF�      PPG �      3
P�      adin�      Spot�      , Pa�      
TX�      oduc�      ug\s�      OFT"�      LOAD�      \spo�      eqio�      #1
�      prod�      plug�      "WEL�      XPLO�      ct\s�      sweq�      " #1�      D pr�      otpl�      u "C�      
TXP�      duct�      g\sw�      HK" �      OAD �      spot�      onf �      1
T�      rodu�      lug\�      APFI�      PLOA�      t\sp�      ftpg�       #1�       pro�      tplu�       "TP�      TXPL�      uct\�      \sws�      I" #�      AD p�      potp�      uf "�      
TX�      oduc�      ug\e�      OT" �      OAD �      spot�      dvf �      1
T�      rodu�      lug\�      K934�      PLOA�      t\sp�      tk94�       #1�       pro�      tplu�       "K9�      TXPL�      uct\�      \atk  H552      XPLOH552      potpH552      K946H552      D prH552      ug\aH552       #1H552      ductH552      k953H552      TXPLH552      spotH552      "K95H552      AD pH552      lug\H552      " #1H552      oducH552      tk96H552      
TXPH552      \spoH552       "SCH552      OAD H552      plugH552      P" #H552      roduH552      sweqH552      LOADH552      tpluH552      c
PH552      ct\sH552      in.pH552      roduH552      swweH552      LOADH552      tpluH552      
PCVH552      \spoH552      tl.pH552      roduH552      swutH552      OAD H552      plugH552      
PCVH552      \spoH552      ld.pH552      roduH552      swprH552      LOADH552      tpluH552      c
PH552      ct\sH552      homeH552       proH552      g\ffH552      CVLOH552      potpH552      .pcH552      ductH552      axtdH552      AD pH552      lug\H552      
PCVH552      \spoH552      sk.pH552      roduH552      swaxH552      LOADH552      tpluH552      c
PH552      ct\sH552      tsk4H552       proH552      g\swH552      CVLOH552      potpH552      .pcH552      ductH552       #�H552      \tptH552      1
TH552      ct\hH552      CFGMH552      D prH552      ftptH552      
TXPH552      \h51H552      AR" H552      prodH552      nrg H552      XPLOH552      510\H552      " #1H552      oducH552      o "MH552      LOADH552      0\sfH552      #1
H552      uct\H552      "MNIH552      AD pH552      sfmnH552      
TXH552      t\h5H552      NJP"H552       proH552      mnmsH552      TXPLH552      h510H552      L" #H552      roduH552      st "H552      PLOAH552      10\sH552       #1H552      ductH552       "TPH552      OAD H552      \sftH552      1
TH552      ct\hH552      TPDAH552      D prH552      psysH552      TXPLH552      h510H552      F" #H552      roduH552      rl "H552      PLOAH552      10\tH552       #1H552      ductH552       "FRH552      OAD H552      \tpfH552      1
TH552      ct\hH552      ORDEH552      D prH552      persH552      
TXPH552      \h51H552      RS" H552      prodH552      fty H552      XPLOH552      510\H552      " #1H552      oducH552      s "TH552      LOADH552      0\tpH552      #1
H552      uct\H552      "CLCH552      AD pH552      tpscH552      
TXH552      t\h5H552      PMA"H552       proH552      smstH552      TXPLH552      h510H552      R" #H552      roduH552      lm "H552      PLOAH552      10\tH552       #1H552      ductH552       "TPH552      OAD H552      \tpdH552      1
TH552      ct\hH552      GRDTH552      D pr           prbd           
TXP           \h51           DT"            prod           odt            XPLO           510\           " #1           oduc           r "T           LOAD           0\sf           #1
           uct\           "SLC           AD p           tpfi           
TXP           \h51           EM"            prod           emd            XPLO           510\           " #1           oduc           r "T             �                         ess            t I)           prod           asde            ! r            usi           rsal           !
I            R83           adin           ersa            Par           OAD            \srg           F  !           
! s           Serv           IF O�          37 R�          Load�          rvo �          I) "�          oduc�          def.�           srv�          ! mi�          IG C�          RDER�          837 �          37
�          ng M�          E, P�          VLOA�          gcor�          PCVL�          migc�          
IF�          R837�          
PCV�          \mig�          f.sv�          LOAD�          core�          NDIF�          fd
�           - M�          ive �          ORDE�          R691�          PRIN�          701 �          ptiv�           I) �          rodu�          pdef�          ! j7�          j703�          E Of�          ORDE�          R691�          PRIN�          703 �          set,�          PCVL�          j703�          NDIF�          
!
�          MIG �          idnc�          ER J�          1 R6�          NT "�           (MI�          void�           "
�          uct\�          f.sv�          706.�          g.fd�          Jog�           R52�          adin�          ched�          ) "�          duct�          f.sv�          jog.�          link�          k I/�          ER J�          7 J5�          
PR�           J85�          /O, �          CVLO�          rcli�          v
E�          ink.�          pprx�          Prox�          ER J�          7 J5�           J68�          adin�           Pro�          "
P�          ct\s�          def.�           smt�          
! a�          Simp�          te
�          R609�           "Lo�          Simp�          te, �          CVLO�          utot�          sv
�          otch�          sths�          AST�           HST�          R794�          ding�          TAST�          
PCV�          \tas�          ���           Ang�          "
P�          ct\t�          sv
�          g.fd�          cp.f�          CP
�          R581�           "Lo�          Modb�           I) �          rodu�          btsv�          F  !�          
!
�          PROF�          
IF �          PRIN�          930 �          O, P�          VLOA�          30\p�          NDIF�          
!
�          FSW �          !
I�          
PR�           J96�          amin�          
PC�          t\j9�          
EN�          fd
�           - T�          Comp�          ER J�          Load�          ol T�          , Pa�          LOAD�          8\gf�          DIF �          !
!�          RCal�          ster�          R J9�          NT "�           (iR�          VMas�           "
�          uct\�          .sv�          92.f�          .fd �          ceNe�          ORDE�          T "L�          (Nad�           WC,�          PCVL�          ndnw�          
END�          d
!�          - La�          I/F�           J59�          adin�          r we�          art �          D pr�          lide�           ! j�           cma�          n ap�          
IF�          J590�          ding�          n ap�          art �          D pr�          pcde�           ! c�           j69�          Torc�          ER J�          Load�          rvoT�          ) "�          duct�          .sv�          CR H�          C H5�          LOAD�          1\sv�          NDIF�          691.�          2.fd�          h fo�          IF O�          RINT�          82 (�          or A�          ) "�          duct�          .sv�          CR H�          C H5�          LOAD�          2\sv�          NDIF�          982.�          0.fd�          h fo�          IF O�          RINT�          80 (�          or S�          ) "�          duct�          .sv�          CR H�          C H5�          LOAD�          0\sv�          NDIF�          580.�          1.fd�           pan�          �j �          !
I�           H54�          T "L�          (Wea�          ) "�          duct�          sv
�          4.fd�          fd -�          C
!�          804�          ing �          us P�          "
P�          ct\j�          sv
�          4.fd�          fd -�          on V�          ORDE�          
PRI�          J996�          ion �          I) "�          oduc�          ef.s�          j996�          mo.f�           Mod�           ORD�          
PR�           R73�          Modi�          ) "�          duct�          .sv�          mo.f�          .fd �          ion�           R65�          H573�          806 �          RINT�          54 (�          n, P�          VLOA�          cz\c�          NDIF  STD   
!
LANG  d - LANG  ol CSTD   
IFSTD   671STD   LoadSTD    (SeSTD    ChaSTD   t I)STD   OAD STD   j671STD   .svSTD   ! j6STD   
! STD   - SeSTD    ChaSTD   IF OSTD   C J6STD   J671STD   RINTSTD   g SVSTD   o HaSTD   e, PSTD   
PCSTD   oducSTD   hdefSTD   IF  STD   d
!STD   .fd STD    funSTD   
IFSTD   683STD   LoadSTD    (StSTD   ctioSTD   I) "STD   D prSTD   83\sSTD   v
ESTD   j683STD   ! j8STD   CD jSTD   utpuSTD    ORDSTD   J619STD   69
STD   oadiSTD   (CD STD   outpSTD    I) STD   AD pSTD   846\STD   sv
STD    j84STD   
! jSTD    M90STD   HiOpSTD    ORDSTD   
PRISTD   ing STD   00iASTD   pt, STD   "
PSTD   roduSTD   m94lSTD   PCVLSTD   uct\STD   idefSTD   IF  STD   d
!STD   .fd STD   InteSTD   
IFSTD   758STD   LoadSTD    (FiSTD   rfacSTD   I) "STD   D prSTD   58\fSTD   sv
STD    j75STD   
! jSTD    FL-STD   IF OSTD   9 J5STD   
PRISTD   ing STD   -netSTD   ) "RBT    proRBT   9\flRBT   v
ERBT   j759OPTN  ! j5OPTN  SafeOPTN  by FOPTN  
IFOPTN  586 OPTN  6
POPTN  adinOPTN  SafeOPTN  by FOPTN  art OPTN  VLOAOPTN  t\j5OPTN  ef.sOPTN  �r4OPTN  IF  OPTN  d
!OPTN  .fd OPTN   TriOPTN  
IF OPTN  25 HOPTN  
PROPTN  dingOPTN  otioOPTN  r, POPTN  
PCOPTN  oducOPTN  gdefOPTN  ORDEOPTN  558OPTN  CVLOOPTN  ct\jOPTN  def.OPTN  F
EOPTN  j625OPTN  ! maOPTN  - PoOPTN  nap OPTN  
IFOPTN  596OPTN  LoadOPTN   (PoOPTN  nap OPTN  art OPTN  VLOAOPTN  t\maOPTN  ef.sDPND    ! DPND  d
!DPND  .fd DPND  PlugDPND  IF ODPND  7
PDPND  adinDPND  PainDPND  n, PDPND  
PCDPND  oducDPND  pdefDPND  IF  DPND  d
!DPND  .fd DPND  tionDPND  I
!DPND  ER RDPND  NT "DPND  R754DPND  tionDPND  I, PDPND  
PCDPND  oducDPND  bskdDPND  NDIFDPND  .fdDPND  12.fDPND  sionDPND  ts
DPND  DER DPND  INT DPND   J91DPND  ion DPND  s, PDPND  
PCCUST  oducCUST  itpdCUST  NDIFCUST  .fdCUST  sdmeCUST  Sys CUST  
!CUST  R SMCUST  J737CUST  RINTCUST  g SMCUST  Dsn CUST  rt ICUST  LOADCUST  \sysCUST  sdsnCUST  NDIFCUST  menuCUST  ! j7CUST  DataCUST  etw.CUST  
IFCUST  740CUST  LoadCUST   (DaCUST  .betCUST   ParCUST  PCVLCUST  uct\CUST  rdefCUST  IF  CUST  d
!CUST  in.fCUST  i UpCUST  
IF CUST  07 HCUST   R72CUST  796 CUST  4 R8CUST  R775CUST  "LoaCUST  7 (ACUST  oad,CUST   "
CUST  prodCUST  in\aCUST  v
ECUST  ascb�      
! �      - TO�      rt
�      DER �      7 R5�      R617�      01 R�       R67�      609 �      INT �       TQS�      oftp�      t I)�      OAD �      tqsp�      v
E�      tqsp�      ! cn�      Cont�      nter�      
IF �      56 J�      NT "�      J756�      lNet�      ce, �      "
P�      rodu�      cnsv�      ENDI�      t.fd�      bdrv�      ther�      iver�      ORDE�      555 �      5 R6�      J757�      58 R�       J59�      688 �      INT �       MOB�      rboa�      r, P�      
PC�      oduc�      mbsv�      ENDI�      rv.f�      h848�      20iA�      
IF �      48
�      oadi�        ���         �      H612�      "Loa�      2 (R�      250F�      ) "�       pro�      2\st�      
EN�      612.�       h61�      -200�      
!�      R H6�      T "L�      613 �      B/18�       I) �      AD p�      613\�      sv
�       h61�      
! e�      EGD �       I/O�      ORDE�      793�      Load�       (EG�      et I�       I) �      AD p�      gd\g�      v
E�      egd.�       cyc�       Cyc�      Trac�      
IF �      22 R�      
PR�      ding�      ycle�      acki�       I) �      AD p�      ycti�      f.sv�       ! c�      
!�      .fd �      hern�      ts
�      DER �      4 H5�      CVTP�      KL J�       PHS�      759 �      1 R6�      J909�      30 J�       J91�      946 �      M R7�      R672�      93 C�        �      $CLA�      ����       ��$�      Z  �      �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          99     ����$FEAT_DEMO U������   �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                            �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �            �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �                �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �$FEAT_DEMOIN         ��   �$FEAT_INDEX         ��   ��$FILECOMP V�������        �$FILESETUP2 W�������  �  N   N �$FILE_AP2BCK 1X������  �)MAKRO900.TP                               %MAKRO900                                 %MAKRO900                                  )MAKRO910.TP                               %MAKRO910                                 %MAKRO910                                  )MAKRO920.TP                               %MAKRO920                                 %MAKRO920                                  )MAKRO930.TP                               %MAKRO930                                 %MAKRO930                                  )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_APPBCK 1X������ 2 �)*.VR                                      %*                                         %                                           )*.PC                                      %FR6:*.PC                                 %                                           )*.TX                                      %FR6:*.TX                                 %                                           )*.FVR                                     %	FR6:*.FVR                                %                                           )*.STM .STM                                %FR:*.STM .STM                            %iPendant Panel                            )*.HTM                                     %FR:*.HTM                                 %                                           )*.GIF                                     %FR:*.GIF                                 %                                           )*.JPG                                     %FR:*.JPG                                 %                                           )*.JS                                      %FR:*.JS                                  %
JavaScript                                )*.CSS                                     %FR:*.CSS                                 %Cascading Style Sheets                    )
ARGNAME.DT                                %FR:\ARGNAME.DT                           %ARGNAME                                   )	PANEL1.DT                                 %FR:PANEL1.DT                             %iPendant Panel                            )	PANEL2.DT                                 %FR:PANEL2.DT                             %iPendant Panel                            )	PANEL3.DT                                 %FR:PANEL3.DT                             %iPendant Panel                            )	PANEL4.DT                                 %FR:PANEL4.DT                             %iPendant Panel                            )SHELL.VR                                  %SHELL                                     %�                                          )ZG_MENUE.VR                               %ZG_MENUE                                  %�                                          )
EINGABE.VR                                %EINGABE                                   %�                                          )SUMM_VAG.DG                               %FR:SUMM_VAG.DG                           %�                                          )TPE_STAT.VR                               %TPE_STAT                                  %�                                          )
TPEINS.XML                                %FR:\TPEINS.XML                           %Custom Toolbar                            )PASSWORD.DT                               %FRS:\PASSWORD.DT                         %Password Config                           )VAGCONF1.XML                              %FR:\VAGCONF1.XML                         %�                                          )EXTSERVO.VR                               %EXTSERVO                                  %�                                          )	IO_SET.DT                                 %FR:\IO_SET.DT                            %�                                          )VWEMZROU.VR                               %VWEMZROU                                  %�                                          )VAGBCKUP.VR                               %VAGBCKUP                                  %�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_DGBCK 1X������ ( �)
SUMMARY.DG                                %MD:SUMMARY.DG                            %Diag Summary                              )
CONSLOG.DG                                %MD:CONSLOG.DG                            %Console log                               )	TPACCN.DG                                 %	TPACCN.DG                                %TP Accounting                             )FR6:IPKDMP.ZIP                            %
IPKDMP.ZIP                               %TP Exception                              )MD:MEMCHECK.DG                            %MD:SUMMARY.DG                            %Memory Data                            �)MD:SHADOW.DG                              %MD:SUMMARY.DG                            %Shadow Changes                        �y�)	FTPLOG.DG                                 %MD:SUMMARY.DG                           %Comment TBD                           \+�)ETHERNET.DG                               %MD:ETHERNET.DG                           %Ethernet Configuration                    )MD:DCSVRFY.DG                             %MD:SUMMARY.DG                           %DCS verify all                        ���)MD:DCSDIFF.DG                             %MD:SUMMARY.DG                           %DCS verify diff                       ���)MD:DCSCHGD1.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �a�)MD:DCSCHGD2.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �a�)MD:DCSCHGD3.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �a�)UPDATES.DAT                               %FRS:\UPDATES.DAT                         %Updates List                              )
PSRBWLD.CM                                %FRS:\PSRBWLD.CM                          %PS_ROBOWELD                               )MD:SMTPLOG.DG                             %MD:SUMMARY.DG                            %SMTP/Email diag                       �@l)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_FRSPRT  �������    �$FILE_MDONLY 1X������    
 �)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_VISBCK 1X������ 
 �)*.VD                                      %FR:\VISION\DATA\*.VD                     %Vision VD file                            )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FMR2_GRP 1Y������� �C4  B�   	                             	 E�� E�@ E�@ E�� E�� E��              	 OHcGPPL�uSL�uSK�y
             	 ?�  ?�  ?�  ?�  ?�  ?�               	 :G:�:G:�:G:�9{��9{��9{��             	 A�  A�  A�  A�  A�  A�  A�  A�  A�  BH   	 C��NC��NC��NB�ƈB�ƈB�ƈ                	                                      	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	 >t�>S��=�h=���>�=��;             	 :�B:{eg:�sX:+N:I9��             	                                      	                                      	 E�  F,D F,D E(p E(p D�               	 ED  E�� E�� D�� D�� DD              C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FMR_CFG Z������� T                                                                                    �$FNO �������F173328               �$FRM_CHKTYP  ����   ������$FROMCHK_MIN        ���  X�$FSSB_CFG [������                                                                           �$FTP_DEF_OW         �    �$FTP_DIRCOMP         �    �$FUNC_SETUP  �������                                                                                  �$GENOVRD_DO        �   �    �$GENOVRD_THR         d   �   d�$GENOV_ENB         �   �$GRAVC_GRP 1\������  �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            ��$GROUP 1b�������                       8�?�              ?�              ?�                  8��q�2ϑf��  ���n��  �ϑc��  4��3q�C�H�l�3DY�    C�  C>                                                             C                 B�                                                                 8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   81�?�              ?�              ?�                  81�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  C�  C�                                                              �                  B�                                             �$GRSMT_GRP 1c�������      C�      C�      C�      C�  �$HOSTC_CFG 1d������ ��                  	FTP       �            �                          172.26.26.230                e                                                                                                       e�                                                                                                      172.26.26.230         e	cfg_fanuc                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �$HOSTENT 1e�������  P!�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !QUICC0                                  !172.26.26.87                      !QUICC1                                  !�                                  !QUICC2                                  !�                                  !ROUTER                                  !172.26.26.1                       !PCJOG                                   !192.168.0.100                     !CAMPRT                                  !192.168.1.10                      !CAMRTR                                  !192.168.1.10                      �$HOSTNAME !�������!KJLTVL111180R01RS--KU1            �$HOSTS_CFG 1d������ �Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                                     	SM                     �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                            �    �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �$HOST_ERR f�������                    �$HOST_PDUSIZ     ^  ��  >�$HOST_PWRD ?������   �  backup        guest         guest         guest         guest         guest         guest         guest         �$HSCDMNGRP 2g������� �      d               K       	P01.05 8   	   	�  �  	�  ]  N  �             	 ���y���2������������             	   	�  �  	�  �  P  <             	 ���y���2���9���V�������             	   �  
�  �  P  �  
�             	 ���j���(���S���������U             	   �  �  �  �  9  �               d 	   	�  �  	�  ]  N  �             	 ���y���2������������                  d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                     �$HSCD_GROUP 2h������      	HSCD01.01         �                  �                  �              �$HSCD_QUPD         �   �$HSCD_UPDTYP  �������   �$HTTP_AUTH 1i�������  <!iPendant                          �                    !KAREL:*                           �                    !KCL:*                             �                    !VISION SETUP                      �                    !�                                  �                    !�                                  �                    !�                                  �                    !�                                  �                    �$HTTP_CTRL j�������                 
 <RFFF9E3                       FRS:DEFAULT               FANUC Web Server             
�$HTTP_PWRD ?������   �  �              �              �              �              �              �              �              �              �$HWR_CONFIG k�������  f                    �$IBGN_CFG l�������       2   @   <#�
<#�
<#�
BH  <#�
<#�
<#�
CH            4   <#�
        �$IBGN_DEV       ���   �$IBGN_ERRIO m�������                �$IBGN_EXDAT n������   �            �$IBGN_EXFLG            �    �$IBGN_FIL o�������                    �$IBGN_FTP p�������                    �  �	MERCATOR  	RECORD    	R_ACHS    	R_ISTW    IBGN  IBG   	SENSPS    TXT   999   	Keine 0                                     %IBSCRECS                               8�%IBSCRECE                               ��           �$IBGN_LMTN  �������                                                                                                                         �$IBGN_SBADR      ���   ��^�x�$IDL_CPU_PCT      B�   BZA��$IDL_MIN_PCT      B�   =��n�$IGNR_IOERR        ���   �$INPT_SIM_DO        ��    �$INTPMODNTOL         ��    �$INTP_PRTY        ��    �$IOLNK 1q�������                                                                                                                                  �$IOMASTER         �    �$IOSLAVE r�������    �$IO_AUTO_CFG         �    �$IO_AUTO_UOP         �    �$IO_CYCLE         �    �$IO_DEF_ASG 1s�������              d                     d                �   c                �   c                  
   c                  
   c                                                                                                                                                                                                                                                                                                                                                                                                                 �$IO_DEF_NUM     ����   �$IO_IPCHE         �   �$IO_RTRY_CNT      ����    �$IO_SCRN_UPD        ��    �$IO_UOP_CFG t�������    �������������������������$ISDT_ISOLC  �������                  �$J23_DSP_ENB  �����������$JOBPROC_ENB         �    �$JOG_GROUP 1u������� 8   d8�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8!�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d81�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8A�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                �$JOG_IN_AUTO      ����    �$JPOSREC_ENB         �    �$KANJI_MASK        ���    �$KAREL_CFG v�������          �$KAREL_ENB         �   �$KCL_LIN_NUM         �   �$KEYLOGGING  ����   d�   �$LANGUAGE �������ENGLISH       �$LGCFG w�������         ��   x  �  �  H  �   '0           �                     MC:\RSCH\00\                 �$LN_DISP x�������                                                    �$LOCTOL      Dz  �A   �$LOGBOOK y�������   d               d  X                                                                                                                                              	LOGBOOK            ��                                                �$LOG_BUFF 1z�������                    d                         d                                                                                                                                                                                                                                                                                                                                                                                   �$LOG_DCS |�������    =���                                        �������������������������������������������������������������$LOG_DIO 1}�������  ������������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ����������������������$LOG_ER_ITM  ������� d                                                                                                                                                                                                                                                                                                                                                                                                                 �$LOG_ER_SEV  �������   �$LOG_ER_TYP  �������                                                                                  �$LOG_REC_RST         �   �$LOG_SCRN_FL 1~�������    �                                                                                                                                                           �$LOG_TPKEY  �������                 �$LONGNAM_ENB         �   �$LUPS_DIGIT         �   �$LU_LOADPROG %�������%UP024                                 �$MAXUALRMNUM       ��   
�$MAX_DIG_PRT        �   �$MCSP ������                                d                �$MCSP_GRP 2�������  �   2     	   �  +  �                         	                                      	                                             	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                     �$MD_LDXDISAB  �����������$MEMO_APNAME ?������� 
 �              �              �              �              �              �              �              �              �              �              �$MISC 1��������  � 	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                         �$MISC_MSTR ��������    �$MISC_SCD 1�������� 
 � 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$MKCFG ��������                       �$MLTARM_CFG �������          �����������������������������$MLT_GRP_DO ��������         ��L��                                                                                                                                        �$MMETPU       ���    �$MNDSP_CMNT         �    �$MNDSP_MST ��������                                              �$MNDSP_POSCF         �   �$MNDSP_PRPMT         �   �$MNDSP_PSTOL 1��������  4@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�$MNSING_CHK         �    �$MODAQ_CFG ��������                             �$MODAQ_DEV 	�������	MC:       �$MODAQ_HSIZE  �������   ��$MODAQ_TASK %�������%$123456789 123456789 123456789 123456  �$MODAQ_TRIG 1��������  l������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ����������$MODAQ_TYPE      ����   �$MODEM_INF 1������� `)AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          �$MONITOR_MSG ?	�������   	EXEC1     	EXEC2     	EXEC3     	EXEC4     	EXEC5     	EXEC6     	EXEC7     	EXEC8     	EXEC9     	EXEC10    	EXEC11    	EXEC12    	EXEC13    	EXEC14    	EXEC15    	EXEC16    	EXEC17    	EXEC18    	EXEC19    	EXEC20    	EXEC21    	EXEC22    	EXEC23    	EXEC24    	EXEC25    	EXEC26    	EXEC27    	EXEC28    	EXEC29    	EXEC30    	EXEC31    	EXEC32    �$MOR_GRP_SV 1�������  ( 	 =���
�?
h=��뿽�/?�;�             	 B�                                  	 B�                                  	                                     �$MOTASK_DATA  �������    �$MPL_NAME !�������!Default Personality (from FD)     �$MRR2_GRP 1����  	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                              �\  �  ��  ��  A�  B  BT  B�   
   �H  ��  ��  A�  B  Bp  B�  C   C   P Dz  E;� E@ D�� D�� D�� C�  C�  Dz      D�� D�� Dz  C�  C�  C�  Dz  D�� C�  E@ D�  D�� D�� Dz  Dz  C�  D�� E;� E;� E@ E/  D�� Dz  C�  C�  E;� D�� E@ E/  E@ D�@ C�  C�  D�� D�  D�� D�  E@ D�� C�  D�� C�  D�� D�  E	� D�  D�� C�  E@ C�  C�  C�  DԀ E@ C�  C�  C�  C�  D�� C�  C�  Dz  C�  C�  C�  D�� E@ C�  C�  C�   P     D�  E;� EZ� E@ E;� EZ� E;�     Dz  E;� EZ� E�� Ez  EZ� E;�     Dz  E;� EZ� EZ� Ez  EZ� E;� D�@ Dz  D�  E�� E;� E�� E�� EZ� E@ D�� E�� E�� EZ� E�  E�  EZ� E@ D�  E�� E�� Ez  Ez  E;� EZ� D�  E@ E�� E�� Ez  Ez  Ez  Ez  E;� E@ E�� E�� E�� Ez  Ez  Ez  E;� E;� E�� E�� E�� Ez  Ez  Ez  E;� E;� E�� E�� E�� Ez  Ez  EZ�  P E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E;� E� E� E� E� E� E� E� EZ� E� E� E� E� E� E� E� Ez  E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E�   DC�*D�+�E�       	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$MRR_GRP 1�������  `     � �     � @D�  D�  ?�  ?�   �?   ?�      @T;gD�  D�                             ;�	l?�   	 ����X�    	 �X^ �,X � � � 	 K��K��eK���K~o�K{GK�M             	                      	   �  �  �  �  �  �  �  �  � 	 ?�;g?��?�;g@
�@
�@T;g                     	 �Iۿ�
��}v�����X���             	 �4  �p  �
=ô  ��  ô               	     >�L����    ���                 	                      �   �   � 	                                 	   ,    �  �  �  M  �  �  � 	                                      	  	'� �  �  I� �  ��             	 :�È:�È:�È:�È:�È:�È=���=���=��� 	  @ @ @ @ @ @             	   �  �  �  �  �  �              �    	                                	   ��  ��  ��  ��  ��  ��  ��  ��  �� 	 @I�?��@�t�@��@�X@��             	 C4  B�  Cf  C�  B�  C�                  ��CR   	  � ���        	        � � H       	 B�  B�  B�  B   B   B                 @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  �� �x @            �   � :              �   ?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  ?      �?            	  (   (   (   P   P   P            	             �>�33       	 ;��;aʤ;r�@;��;�	�<$D             	                       A0              ?�   �    ?@    ?fff?@  ?&ff?    	 A�A�A�@�,@�,@�,            CR    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	     D�� E��     E9� E�0              	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 G=�GW�G�QFcNfC��AFBC           	                                                                                       Ap  �?��                    �p  BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                      	                                      	     ?��                             	                                      	             Ġ      �k               	 C�  D�` Ca                           	 ?��    ���?�ؿ��@I�             	 C��CHf�CW�FB�1B-v�=���             	 É����XR���u                     	 �ę����AP��Blz��X��                 	 ¡�R�d�
Ák�BU(���  ��              	 K���JGp@KÌH�� I%K�AP               	 L)-yL!�GKӕ#HP� H�R�AP               	 L(�L&��J�3$H㞀H���A�               	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	     G�?                              	     C�?�                             	     Ć�                             	     CV��                             	                                      	 �                                   	                                      	                                      	 ( 	 �`��                    ��������� 	     �1V                ��������� 	         3>�            ��������� 	             3��v        ��������� 	             ��v3�g�    ��������� 	             �!�;�%D93ҵ���������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	       �                             	                                      	                �                     	               8  t                 	                                      	                                      	                                      	 ( 	                             	                             	      �                      	                             	            O�                	            �e 3�             	                             	                             	                                 2 D�         Ep         E�         B�  A   A�  C�  D  A   @�                                      �                                               D� D�         �                                            D�         Ep         E�                                                                                     ?�  ?�              	                                
                                                                                                                                                                                                                                                                                          	     ��            �̿��      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 C_ff                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C��                                          	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 CU��                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$MSKCFMAP  �������                               �$MSKCONREL         �   �$MSKEXCFENB         
�    �$MSKEXCFFNC         
�   �$MSKJOGOVLIM         d�   d�$MSKKEY         �   �$MSKKEY_PANL             �$MSKRUNOVLIM         �   �$MSKSFSPDTYP         
�    �$MSKSIGN         �   �$MSKT1MOTLIM         d�   �$MSK_CE_GRP 1��������  \     	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                        �$MSQZ_EDIT      ����    �$MTCOM_CFG 1��������         
       
       
       
       
       
       
       
�$MT_ARC_ENB         �   �$MUAP_CPLENB         �    �$NOCHECK ?�������  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �$NO_WAIT_LN        ���   �$NUM_RSPACE  �������     
   
   
   
   
   
   
   
�$ODRDSP_ENB         �    �$OFFSET_CART         �    �$OFFSET_DIS         �    �$OPEN_FILES     
   ��   
�$OPTION_IO         �   �$OPTM_PRG %�������%$************************************  �$OPWORK ��������    �� �� ��       ���                        	 �                      �      ��$ORG_DSBL  �������                                  �$ORIENTTOL      C�  �A   �$OUT_SIM_DO        �    �$OVRDSLCT ��������    ������   
   
   
   
    �$OVRD_PEXE         �    �$OVRD_RATE         d�   �$OVRD_SETUP ��������     
 ����������������������������������������     
 �����������������������������������������$PARAM2_GRP 1���� 	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                              �\  �  ��  ��  A�  B  BT  B�   
   �H  ��  ��  A�  B  Bp  B�  C   C   P Dz  E;� E@ D�� D�� D�� C�  C�  Dz      D�� D�� Dz  C�  C�  C�  Dz  D�� C�  E@ D�  D�� D�� Dz  Dz  C�  D�� E;� E;� E@ E/  D�� Dz  C�  C�  E;� D�� E@ E/  E@ D�@ C�  C�  D�� D�  D�� D�  E@ D�� C�  D�� C�  D�� D�  E	� D�  D�� C�  E@ C�  C�  C�  DԀ E@ C�  C�  C�  C�  D�� C�  C�  Dz  C�  C�  C�  D�� E@ C�  C�  C�   P     D�  E;� EZ� E@ E;� EZ� E;�     Dz  E;� EZ� E�� Ez  EZ� E;�     Dz  E;� EZ� EZ� Ez  EZ� E;� D�@ Dz  D�  E�� E;� E�� E�� EZ� E@ D�� E�� E�� EZ� E�  E�  EZ� E@ D�  E�� E�� Ez  Ez  E;� EZ� D�  E@ E�� E�� Ez  Ez  Ez  Ez  E;� E@ E�� E�� E�� Ez  Ez  Ez  E;� E;� E�� E�� E�� Ez  Ez  Ez  E;� E;� E�� E�� E�� Ez  Ez  EZ�  P E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E;� E� E� E� E� E� E� E� EZ� E� E� E� E� E� E� E� Ez  E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E� E�                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$PARAM_GROUP 1�gX�� `     � �     � @D�  D�  ?�  ?�   �?   ?�      C>  D�  D�                             ;�	l?�   	 ����X�    	 �X^ �,X � � � 	 H��H�ffH�  H��H�WH-��             	                      	   �  �  �  �  �  �  �  �  � 	 B�  B�  B�  B�  B�  C>                       	 �4  �p  �
=ô  ��  ô               	 �4  �p  �
=ô  ��  ô               	     A�8�¼r�    «�C                 	                      �   �   � 	                                 	   ,    �  �  �  M  �  �  � 	                                      	  	'� �  �  I� �  ��             	 =���=���=���=���=���=���=���=���=��� 	  @ @ @ @ @ @             	   �  �  �  �  �  �              �    	                                	   ��  ��  ��  ��  ��  ��  ��  ��  �� 	 C4  B�  Cf  C�  B�  C�               	 C4  B�  Cf  C�  B�  C�                  ��CR   	       ��        	        � � H       	 B�  B�  B�  B   B   B                 @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  �� �x @            �   � :             �   ?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  ?      �?            	  (   (   (   P   P   P            	             �>�33       	 ;��;aʤ;r�@;��;�	�<$D             	                       A0              ?�   �    ?@    ?fff?@  ?&ff?    	 A�A�A�@�,@�,@�,            CR    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	     D�� E��     E9� E�0              	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                       Ap  �?��                    �p  BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                      	                                      	     ?��                             	                                      	             Ġ      �k               	 C�  D�` Ca                           	 ?��    ���?�ؿ��@I�             	 C��CHf�CW�FB�1B-v�=���             	 É����XR���u                     	 �ę����AP��Blz��X��                 	 ¡�R�d�
Ák�BU(���  ��              	 K���JGp@KÌH�� I%K�AP               	 L)-yL!�GKӕ#HP� H�R�AP               	 L(�L&��J�3$H㞀H���A�               	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	     G�?                              	     C�?�                             	     Ć�                             	     CV��                             	                                      	 �                                   	                                      	                                      	 ( 	 �`��                    ��������� 	     �1V                ��������� 	         3>�            ��������� 	             3��v        ��������� 	             ��v3�g�    ��������� 	             �!�;�%D93ҵ���������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	       �                             	                                      	                �                     	               8  t                 	                                      	                                      	                                      	 ( 	                             	                             	      �                      	                             	            O�                	            �e 3�             	                             	                             	                                 2 D�         Ep         E�         B�  A   A�  C�  D  A   @�                                                                                      D� D�                                                                                                                                                                      ?�  ?�              	                                
                                                                                                                                                                                                                                                                                          	     ��            �̿��      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 C_ff                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C��                                          	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 CU��                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$PARAM_MENU ?�������  DEFPULSE              	WAITTMOUT             RCVTMOUT              SHELL_WRK.$CUR_STYLE  SHELL_WRK.$CUR_OPTA   SHELL_WRK.$CUR_OPTB   SHELL_WRK.$CUR_OPTC   SHELL_WRK.$CUR_DECSN  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PASSREL_ID      ���   �    �$PAUSE_PROG %�������%�                                      �$PCCRT         �    �$PCCRT_HOST !�������!PCCRT                             �$PCTP         �    �$PCTP_HOST !�������!PCTP                              �$PC_TIMEOUT      ����   �$PGDEBUG  �������    �$PGINP_FLMSK      ����    �$PGINP_FLTR      ����   �$PGINP_PGATR  �������                     �$PGINP_PGCHK      ����   �$PGINP_TYPE ?������  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PGINP_WORD ?	�������  	FOLGE     	UP        	MAKRO     	SUCHL     	MAKROSP   �$PGTRACECTL 1�������� 
    � �   K L   � �   � �                               �$PGTRACEDT Q�������� 
D � 	   	   	   	   	   	   	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  	� c  	� d  	� e  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	� �  	   	 	  	 
     	   	   	   	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	   	   	      	   	   	   	   	   	   	   	   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   	 	  	 
     	               	   	   	    � 	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  �   	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    ��    	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    T   T   T 	  	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   T 
  T   T   T   T   }   }   U   ]   }   �   }   �   �   �   �   �   �   �   �   �   �   �   �   �    �   �   �   �   �   �   �   � 	  � 
  	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /   � � K  � L  � M  � N  � O  � P  � Q  � R  � S  � T  � U  ��    �   �   �   �   �   �   �   �   � 	  � 
  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �    � !  � "  � #  � $  � %  � &  � '  � (  � )  � *  � +  � ,  � -  � .  � /  � 0  � 1  � 2  � 3  � 4  � 5  � 6  � 7  � 8  � 9  � :  � ;  � <  � =  � >  � ?  � @  � A  � B  � C  � D  � E  � F  � G  � H  � I  � J  � K  � L  � M  � N  � O  � P  � Q  � R  � S  � T  � U  ��    �   �   �   �   �   �   �   �   � 	  � 
  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �    � !  � "  � #  � $  � %  � &  � '  � (  � )  � *  � +  � ,  � -  � .  � /  � 0  � 1  � 2  � 3  � 4  � 5  � 6  � 7  � 8  � 9  � :  � ;  � <  � =  � >  � ?  � @  � A  � B  � C  � D  � E  � F  � G  � H  � I  � J  � K  � L  � M  � N  � O  � P  � Q  � R  � S  � T  � U  ��    � ;  � <  � =  � >  � ?  � @  � A  � B  � C  � D  � E  � F  � G  � H  � I  � J   � 	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  ��    	�   	�   	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +  	� ,  	� -  	� .  	� /  	� 0  	� 1  	� 2  	� 3  	� 4  	� 5  	� 6  	� 7  	� 8  	� 9  	� :  	� ;  	� <  	� =  	� >  	� ?  	� @  	� A  	� B  	� C  	� D  	� E  	� F  	� G  	� H  	� I  	� J  	� K  	� L  	� M  	� N  	� O  	� P  	� Q  	� R  	� S  	� T  	� U  	� V  	� W  	� X  	� Y  	� Z  	� [  	� \  	� ]  	� ^  	� _  	� `  	� a  	� b  ��    �   ��    �   ��    	�   	�   	�   	�   	�   	�   	� 	  	� 
  	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�   	�    	� !  	� "  	� #  	� $  	� %  	� &  	� '  	� (  	� )  	� *  	� +   � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    �$PGTRACELEN       ��   ��$PGTRACE_UP ��������   ����$PG_CFG ��������       ����                                                      �$PG_DEFSPD ��������  �     ��$PING_CTRL ��������      8       �$PIPE_CONFIG �����������                   �$PLID_CFG ��������   �$PLID_GRP 1������� �   CH�����    A�  G�G G�7�F�, A�  D	�          �   d      d      d   d   d   d         � 	                                    	                 ´  ´               	                 B�  B�               	                 ´  ´               	                 B�  B�               	                 B��B>�e             	                                      	                 <,1<49X             	                                      	                                      	                                      	                 <,1<49X             	                                      	                                      	                 Dz  Dz                      
 C  @�b���� A��H�x�H�K�G�j                     	                                      	                                      	                                      	                                      	                 >V�>W�             	                                      	                                      	                                        !    
V7.10beta1         @�33@2�\@;�CR    C>  CW  B�    D�� D�� D0�   D�  D�� Dj  C2  A�  B�  CR  C]  Ap     B�  B�  B�ffCX(�B!33BffA�  B\  B\  B,  B\ffB\��B��n�}��v8    ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ����$PLID_KNOW_M         �   �$PLID_SV ���������        
                                                                                  	                                      	                                        d      d   d    �$PLIM_GRP 1��������  lCR   	       ��        	        � � H       �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���$PLMR_GRP 1��������  T        B�  C  CR      C��  
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�              �$PLST_GRP1 1�������� 
 0Vacia             C�N��&����B��H��]H��nG�=Llena             C  @�b���� A��H�x�H�K�G�j�                  CR                          �                  CR                          �                  CR                          �                  CR                          �                  CR                          �                  CR                          �                  CR                          �                  CR                          �$PLST_GRP2 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP3 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP4 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP5 1��������  0�                  �<                         �$PLST_GRP6 1��������  0�                  �<                         �$PLST_GRP7 1��������  0�                  �<                         �$PLST_GRP8 1��������  0�                  �<                         �$PLST_GRPMAD        �   �$PLST_PARNUM  �������                              �$PLST_SCHMAD         �   
�$PLST_SCHNUM         �   
�$PLST_UPDNUM  �������                          �$PLS_CMP_LIM  ����  '�   �$PLS_ER_CHK  ���� ���    �$PLS_ER_LIM  ����  '�   �$PLS_ER_RST         �    �$PL_MOD         �   �$PL_MOD_ST         �   �$PL_RES_G1 1�������� 
                                 C  D8�cD8�cC�>,IB��IB��H%#                                                                                                                                                                                                                                                           �$PL_RES_G2 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G3 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G4 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G5 1��������                                  �$PL_RES_G6 1��������                                  �$PL_RES_G7 1��������                                  �$PL_RES_G8 1��������                                  �$PL_RES_V 1�������   �  �^�`�^h�]�T�]���$PL_THR_INRT         d�   d�$PL_THR_MASS         d�   Z�$PL_THR_MMNT         d�   Z�$PMON_QUEUE ��������       �      �$PM_GRP 2�������  4      A�  @�                    B�           �$PNS_CUR_LIN        ���    �$PNS_END_CUR         �    �$PNS_END_EXE         �    �$PNS_NUMBER        ���    �$PNS_OPTION         �   �$PNS_PROGRAM %�������%PNS                                   �$PNS_TASK_ID        ���    �$POCFG ��������                                      �$PODATA_GRP 1�������� @ �[   # 2  2   " + 0    !   " + 0    !   " + 0    !   " + 0    ! 0    !   " + 0    !  2                                                    �J    2 }}}}} 2     !    " + 0    !    " + 0    !    " + 0    !    " + 0    !    " + 0 2                                                    �J    2 }}}}} 2     !    " + 0    !    " + 0    !    " + 0    !    " + 0    !    " + 0 2                                                    �L    2 }}}}} 2  + 0    !    " + 0    !    " + 0    !    " + 0    !    " + 0    !    " 2                                                   �$POINFO_GRP 1�������� �     �                                                                                                                                                                                                                                                                                                                                                                                                                 �$POIO_GRP 1��������             �$POS_EDIT ��������                               �$POWERFL            �    �$PRGADJ ��������A�  A�  A�  ?   ?   ?      d    �$PRGNS_CFG ��������?�             @   <@�             %�                                                            �$PRGNS_GRP 2�������� �  \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                     �$PRGNS_PREF ��������      
    �$PRIORITY         ��   ��$PRMPDSPON            �    �$PRMPDSPOUT        �   �    �$PRODUCT_ID �������                       �$PROGGRP_TGL      ����    �$PROTOENT 1��������  (!AF_INET                              !tcp                                  !udp                                  !icmp                                 �$PROXY_CFG ��������  �    )� ****************************************   �)� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** �$PRO_CFG ��������    %�                                                          >�%�        ****/**/**/ **:**:**      %�                                         �                        A�    ,  �                                                                                     �$PRO_PREF ��������      
      �$PRPORT_NUM        �   �$PR_CARTREP  �������    �$PSKSTAT         �    �$PSSAVE ��������	2600H601                                              !�                                  !�                                  �                  	�          �        �                         �                      e�                                                                                                      �              !�                                  �$PSSAVE_GRP 1��������    �%��                  ���������������������$PS_CONFIG ��������                     
          �  �   �h+ �$PS_CP_CFG 2��������                                                         �$PS_CP_GRP 2�������   �         U$58���?W?|K;� '?O�>)��?�/?�J���P�pDa�;BjR�D���    8���?W?|K;� '?O�>)��?�/?�J���P�pDa�;BjR�D���        8�?�              ?�              ?�                  q8 n    ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������       �$PS_MOTION 2�������� 
�                                %�                                      %�                                                                                                                  8�?�              ?�              ?�                                                                                                                                                                                                                                                                                                                             ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   EL %�                                    '���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                      %�                                   �%��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   ��%�                                      ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                      %�                                   ~h��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   %�                                      ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   N ]%�                                   �{��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                     %�                                   � ���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   ��%�                                   �
���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   ock%�                                   me=��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$PURGE_ENBL         �   �$PWFENBDO            �    �$PWF_IO        �   �$PWRUP_DELAY ��������       �$PWR_HOT %������   �%�                                      �$PWR_NORMAL %�������%�                                      �$PWR_SEMI %�������%�                                      �$QSKIP_GRP 1��������  x 	                                      	                                                                              	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ����������������������������������������������������������$RBTIF      ����    �$RCVTMOUT        ��  ��$RDCR_GRP 1������� � 	 E�%SE�E�B�D�]�D�W�D��             	 ŏ����J    ċ���94F�{��             	                                      	 ;��;aʤ;r�@;��;�	�<$D                    	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                   �$RDIO_TYPE  �������                                  �$REFPOS1 1�������� 
 x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS2 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS3 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS4 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS5 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS6 1��������  x�                                  	                                      	                                         �$REFPOS7 1��������  x�                                  	                                      	                                         �$REFPOS8 1��������  x�                                  	                                      	                                         �$REFPOSMASK 1��������     
   
   
   
   
   
   
   
�$REFPOSMAXNO  �������     
                     �$REMOTE  �������   �$REMOTE_CFG ��������          �$REPL_RANGE      ����   �$REPOWER ��������    �$RESM_DRYPRG %�������%�                                      �$RESTART ��������            �$RESUME_PROG %�������%�                                      �$RE_EXEC_ENB         �   �$RGSPD_PREXE         �    �$RGTDB_PREXE         �    �$RGTRM_PREXE         �    �$RMT_MASTER  �������    �$ROBOT_ISOLC  �������                 �$ROBOT_NAME �������KJLTVL111180R01       HTML�$ROB_ORD_NUM ?�������  H601 8H895  H895  H895     ���    ��    �|     ��$RPC_TIMEOUT      ����   x�$RS232_CFG 1��������  LTEACH PENDANT                                  �                  Maintenance Conso                          "   �                  	Unbenutzt                                      �                  	Unbenutzt                                      �                  �$RS232_NPORT        �   �$RSCH_LOG ��������       		RSCH          �$RSMAVAILNUM        ��   �$RSPACE1 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                    ���������  ����������                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE2 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE3 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE4 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE5 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE6 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE7 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE8 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACEG ��������                           
 
                                                                                  ������������������������������������������������������������                                                                                                              d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������  `                  @   @   @                                                                           �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                ����������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  ��������������������� 
                                         �$RSPACE_MODE  �������    �$RSPACE_S ��������                                                                                                                          	                                     �$RSPCWORK_AD  ��������@�$RSR  �������                  �$RSR_INTVAL        ��    �$RSR_OPTION         �   �$RTCFG ��������                      ?          �  �   �$RV_DATA_GRP 2�������   � D  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SAF_DO_PULS  ����   �������$SCAN_TIME        ��   �$SCR ����8		      
      
               
                                                                                                                                                                                                                                                                             �         2   2   
   
   d   
   d   2   d                        @                                                                          
                               P       
�� @B     T                                                                                    T D��                                                                                                                                                                                                                                                                                                                                                            @                    




                                             @         ;�o             p              
�t� �Di                     �� �                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                  �                                 0    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                                                                                                                                                                                                  �           �  �  � � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                   T                                                                                                                                                                                                                                                                                                                                                      �                                                       ��                                     	12345678    `!B  �            T                                                                                      T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T BH                                                                                                                                                                                                                                                                                                                                               T ;�j                                                                                                                                                                                                                                                                                                                                             T D�                                                                                                                                                                                                                                                                                                                                               T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   "CH  A�               �          2                   
   d   
  �  	�     2                                                                                                       p  �                                  �                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                                                                                                                                                                                                                                                                                                                                                     �$SCR_GRP 1��� t �            	    � 	    � 	                                  	                                	                                     �      D�` D�                   �     �                            R-2000iB/210F 567890  	R-2000iX  	RB21 678      
V06.10         	          	   
   
   
           	          �       �              	      	          � 	                                                                                                             ��H� 	     	    ��      O�'C��D	��D���Cw�@�a�B�,m 	 @�����AA��	@���©��B�                     >�7C�
D	��D��� 	                                                            	                                         	                      h  �X��     	 B���B�  B�  B�  B�  B�  B�  B�  B�   	 A   A   A   A   A   A   @   @   @    	 @�  @�  @�  @�  @�  @�  ?�  ?�  ?�   	 BH  BH  BH  BH  BH  BH  A   A   A    	 F@ F�` F�`                          	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                            
                                         ?�  @�  @&��                         	 @�  @�  @�  @�  @�  @�  B�  B�  B�  12345678901234567890                                                  A�                	                    	                                                                                                                                           P P P ( ( (                                                        �           	 	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	 B���                                                         	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	 BS��                                                         	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	                                                              	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �$SEL_DEFAULT        ���   �$SEMIPOWERFL         �   �$SEMIPWFDO         �    �$SERVENT 1�������  L!DUM_EIP                             �j!AF_INET                           !FTP                                  !AF_INET                           !�                                    �!AF_INET                           !RPC_MAIN                            �!AF_INET                           !RPC_VISN                            �!AF_INET                           !TP_INPUT                            �d!AF_INET                           !
PMON_PROXY                          �e!AF_INET                           !TP_PROXY                            �f!AF_INET                           !RDM_SRV                             �g!AF_INET                           !R90                                 �h!AF_INET                           !
RPCM_PROXY                          �i!AF_INET                           !RLSYNC                              8!AF_INET                           !ROSIP                               �4!AF_INET                           !
CETP_MTCOM                          �k!AF_INET                           !	CETP_CONS                           �l!AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           �$SERVICE_KL ?%������  (%SVCPRG1                               %SVCPRG2                               %SVCPRG3                               %SVCPRG4                               %SVCPRG5                               %SVCPRG6                               %SVCPRG7                               %SVCPRG8                               %SVCPRG9                               %SVCPRG10                              %SVCPRG11                              %SVCPRG12                              %SVCPRG13                              %SVCPRG14                              %SVCPRG15                              %SVCPRG16                              %SVCPRG17                              %SVCPRG18                              %SVCPRG19                              %SVCPRG20                              %SVCPRG21                              %SVCPRG22                              %SVCPRG23                              %SVCPRG24                              %SVCPRG25                              %SVCPRG26                              %SVCPRG27                              %SVCPRG28                              %SVCPRG29                              %SVCPRG30                              �$SERVICE_PRG ?%������  (%                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       �$SERV_DEV �������MC:           ����$SERV_MAIL      ����    �$SERV_OUTPUT      ����    �$SERV_REC 1�������   �     o 	    #   $   $   %                   	                    	                	                                	                                      
 �W��H6 2    	                         ��������� 	      �   �   �  �  W��������� 	    =   b�������v����  ?��������� 	   �       �  �  v���������W��O6 2    	                         ��������� 	      �   �   �  �  V��������� 	    =   b�������v����  ?��������� 	   ����    �  g  S���������W��[6 2    	                    ��������� 	      �  $   9  j  X��������� 	    =   b�������v����  ?��������� 	 �������F  �  r  �  ����������W��a6 2    	          &          ��������� 	      �  C   2  �  ���������� 	    =   b�������v����  ?��������� 	 ����     |  �  �  $���������W��p6 2    	          /          ��������� 	    	  _  `   -  �  ���������� 	    =   b�������v����  ?��������� 	 �������  �  n  
e  ����������W�J�6 2    	                   ��������� 	       �   #      ��������� 	    9   V�������n����  Q��������� 	 �������   U  ������������������W��u6 2    	                    ��������� 	       �      �   �  w��������� 	 ����   ^����   �����   f��������� 	 �������  2  	u���X  ���������W��.6 2    	    	   $   Q   D   *   6��������� 	    E  \      �  �  ���������� 	 ����   _����   �����   f��������� 	 �������  0  m���?  ]���������W��26 2    	       *   C         ���������� 	    f       �    Q��������� 	    =   b�������v����  ?��������� 	   <���M  �  W  �  	���������W��66 2    	                         ��������� 	      �   �   �  �  u��������� 	    =   b�������v����  ?��������� 	   �����  >  '  �  $���������    
 �W��O6 2    	                         ��������� 	      �   �   �  �  V��������� 	    =   b�������v����  ?��������� 	   ����    �  g  S���������W��p6 2    	          /          ��������� 	    	  _  `   -  �  ���������� 	    =   b�������v����  ?��������� 	 �������  �  n  
e  ����������W��a6 2    	          &          ��������� 	      �  C   2  �  ���������� 	    =   b�������v����  ?��������� 	 ����     |  �  �  $���������W��[6 2    	                    ��������� 	      �  $   9  j  X��������� 	    =   b�������v����  ?��������� 	 �������F  �  r  �  ����������W��H6 2    	                         ��������� 	      �   �   �  �  W��������� 	    =   b�������v����  ?��������� 	   �       �  �  v���������W��66 2    	                         ��������� 	      �   �   �  �  u��������� 	    =   b�������v����  ?��������� 	   �����  >  '  �  $���������W��26 2    	       *   C         ���������� 	    f       �    Q��������� 	    =   b�������v����  ?��������� 	   <���M  �  W  �  	���������W�]z6 2    	                         ��������� 	          �   �  �  ���������� 	    =   b�������w����  =��������� 	    �   j  �  �  �  O���������W��.6 2    	    	   $   Q   D   *   6��������� 	    E  \      �  �  ���������� 	 ����   _����   �����   f��������� 	 �������  0  m���?  ]���������W�]�6 2    	                         ��������� 	          �   �  �  ���������� 	    =   b�������w����  =��������� 	    b   ;  �  k  x  ����������   4 	                                     	                                      	                                     	                                      
 �J���6�     	   ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������K�3�6 2     	   v������������������������ 	     ������������������������ 	   ������������������������� 	     ������������������������N� �6   @  	   ^������������������������ 	     ������������������������ 	   :������������������������ 	     ������������������������REN�6 2     	   ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������RER�6 2     	   ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������W�[�6 2    	   	M������������������������ 	     ������������������������ 	   ������������������������ 	     ��������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������    
 �W��66 2    	     ������������������������ 	     ������������������������ 	   T������������������������ 	     ������������������������W�[�6 2    	    ������������������������� 	     ������������������������ 	   ������������������������ 	     ������������������������W�[�6 2    	     ������������������������ 	     ������������������������ 	   ,������������������������ 	     ������������������������W�[�6 2    	   	M������������������������ 	     ������������������������ 	   ������������������������ 	     ������������������������W�[�6      	     ������������������������ 	     ������������������������ 	   ������������������������� 	     ������������������������W�[�6      	    ������������������������� 	     ������������������������ 	   ������������������������ 	     ������������������������W�[|6 2     	    ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������Iq-k6    	     ������������������������ 	     ������������������������ 	   &������������������������� 	     ������������������������W��6 2    	   ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������K,�6�     	   ������������������������� 	     ������������������������ 	    ������������������������� 	     ������������������������   - 	                                     	                                      	                                     	                                      
 �J.76r _     	   ������������������������� 	     ������������������������ 	   '@������������������������ 	     ������������������������R�&�6    	   ������������������������� 	     ������������������������ 	   R������������������������� 	     ������������������������W�[�6 2    	   .������������������������ 	     ������������������������ 	   'h������������������������ 	     ��������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������    
 �W�[�6 2    	   .������������������������ 	     ������������������������ 	   'h������������������������ 	     ������������������������W�[�6 2    	     ������������������������ 	     ������������������������ 	   'h������������������������ 	     ������������������������W�[�6      	     ������������������������ 	     ������������������������ 	   'm������������������������ 	     ������������������������W�[�6      	   &������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������W�[|6 2     	   &������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������S���6    	   &������������������������ 	     ������������������������ 	   ������������������������� 	     ������������������������W��6 2    	     ������������������������ 	     ������������������������ 	   &������������������������� 	     ��������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     	                                      	                                      	                                      	                                      
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_RV 1�������   �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_TOP10 1�������   � 
 6 2   $6    56 *   6�   6r _   6�   6    6�   6T   6    �$SERV_TYPE      ����    �$SHELL_CFG ��������                                                                %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                                       �  �   %                                                                                                     �         �   2   d                                �$SHELL_CHK 1��������                                                                                                                                                                                                                                                                                                                                                                                  �$SHELL_COMM ��������                        �$SHFTOV_ENB         �    �$SHOW_REG_UI         �    �$SIMWAITENB            �    �$SIMWAITOUT        �   �    �$SIMWAITTIM       ��   �    �$SIMWAITVAL            �    �$SI_UNIT_ENB         �   �$SLC_RETRY         �   �$SMB_HDDN 2��������    ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  �������������������������$SMON_ALIAS ?e������ ( he�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      �$SMON_DEFPRO ������ *SYSTEM*    ��$SMON_RECALL ?}������ ( �}�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              �$SNPX_ASG 1�������� P 0 '%R[1]@1.1                              ?�      %                                    <�Q?�      %                                    _*_?�      %                                    �o�?�      %                                     .�?�      %                                    �� ?�      %                                    ��#?�      %                                    � �?�      %                                    $�E?�      %                                    �K?�      %                                    �8?�      %                                    �0�?�      %                                    !�0?�      %                                     t�?�      %                                    �0?�      %                                    � �?�      %                                    /�?�      %                                    v�?�      %                                    !�2?�      %                                    !̈́?�      %                                    � ?�      %                                    ��?�      %                                     lG?�      %                                    　?�      %                                    Q�?�      %                                    Q<?�      %                                    �� ?�      %                                     ?�      %                                      ?�      %                                    ���?�      %                                     $?�      %                                    &�?�      %                                    2�Y?�      %                                    �ϴ?�      %                                    ?�?�      %                                    ��?�      %                                    � ?�      %                                    �|x?�      %                                    	?�      %                                    n�M?�      %                                    �	�?�      %                                    ��?�      %                                    J�\?�      %                                    �?�      %                                    �?�      %                                    ?5O?�      %                                    O�O?�      %                                    ]o�?�      %                                    v�?�      %                                    zb8?�      %                                    ޒ�?�      %                                    �C?�      %                                    ���?�      %                                     � ?�      %                                    ?�      %                                    ���?�      %                                    �AJ?�      %                                    ��?�      %                                    ��%?�      %                                    �A/?�      %                                    �4�?�      %                                    ~j?�      %                                    @?�      %                                    �I�?�      %                                    �>w?�      %                                    �N�?�      %                                    R�?�      %                                    ���?�      %                                    ��?�      %                                    ���?�      %                                    �6 ?�      %                                    ��?�      %                                     |?�      %                                     '8?�      %                                       ?�      %                                    ��?�      %                                      ?�      %                                       ?�      %                                    �#t?�      %                                    ��\?�  �$SNPX_PARAM ��������  �	�             P                           ��$SOFT_KB_CFG        ���    �$SOPIN_SIM  �������                                                  �$SRVQSTP_DSB  �������                                  �$SSR ������� � & FOLGE011 .......................0006        �$STHI_CHANGE         �    �$STHI_GRPNUM         �    �$STOP_ON_ERR         �    �$STOP_PTN ������C �$STRING_PRM         �   �$SVDT_GRP 1�������    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                   �$SVPRG_COUNT        ��    �$SVPRG_ENB         �    �$SVPRM_ENB         �    �$SVPRM_UPD 1������� T  
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                     �$SV_CTRL_NUM        
�   �$SV_GUN_CTRL 2��������                 /   /   
               4   4   
                        
                           
                           
�$SYSDEBUG  ����   d�    �$SYSDSP_PASS       B?�    �$SYSLOG ��������         �^��                      �       UD1:\SYSLOG               �$SYSLOG_MPC ��������                                    �       UD1:\SYSLOG2              �$SYSLOG_SAV ��������                     UD1:\SYSLOGSV         �$SYSTEM_TIME 1��������  ( @�U     0ȩ        &O�                 @�U     0�        &O�                 @�U     0�        &O�                 @�U     0�        &O�                �$T1SVGUNSPD        '�   ��$TASK_OPTION  ������   �   �$TA_DISP_ENB         �    �$TBCCFG ��������                                                 `                             	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                                                                	                                      	                                      	                                         ��������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������    �$TBCSG_GRP 2��������  �    
 ?͈?͈?͈?͈?͈?͈?͈?͈?͈?͈ 
 ?͈?͈?͈?͈?͈?͈?͈?͈?͈?͈ 
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ��� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������A��*SYSTEM*   V8.2306       4/24/2014 A t  *SYSTEM* *SYSTEM*  F�TBCPARAM_T   �$MC_MAX_TRQ  $MAX_TRQ_MGN  $MC_GRAV_MGN  $MC_STAL_MGN  $MC_BRK_MGN  $MC_NOLD_MGN  $SHORTMO_LIM  $SHORTMO_MGN  $MC_NOLD_TRQ  $J_LIN  $SPL1  $SPL2  $SPL3  $SPL4  $SPL5  $SPL6  $SPL7  $SPL8   ��TBC_GRP_T � $TBC_ACCEL1  $TBC_ACCEL2  $TBC_PATH1  $TBC_PATH2  $PATH_RATIO  $TBC_PARAM 2  	$CNT_SCALE  $SHORTMO_SCL  $MIN_ACC_UCA  $MIN_CAT_UMA  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2L_UPR_ANG  $J2L_LWR_ANG  $J2L_UPR_MGN  $J2L_LWR_MGN  $R_F2LSHRT  $R_F2LLONG  $MIN_F2LSHRT  $MIN_F2LLONG  $MIN_ACRL_S  $MIN_ACRL_L  $MIN_PAYLOAD  $HVAL   $HMGN   $FLEXL   ��TBJ_ACC_T  :$ACC_LEN1  $ACC_LEN2  $DEC_LEN1  $DEC_LEN2  $ACCEL_RATIO  $DECEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $F1DEC_I  $F2DEC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$DECTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT_ACC   	$J_STAT_DEC   	$M_STAT_ACC  $M_STAT_DEC  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $DEC2_STP   $AT_MODE  $AT_AXS   	$AC_ACC   	$AC_DEC   	$JK_ACC   	$JK_DEC   	$VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AA1  $AA2  $AA3  $AA4  $AA5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM  ��TBJCFG_T  � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $UPDATE_TIME  $TBJ_SELECT  $TBJ_STAT   $TJ 2 $JERK_CTRL  $MOTN_INF  $TBJ_DEBUG  $HAND_VB   �TBJOP_GRP_T  $ $F2MGN  $MINF2  $COMP_SW  :�TBPARAM_T � $$MR_MAX_TRQ  $MR_STAL_TRQ  $MR_BRK_TRQ  $MR_BRK_VEL  $MR_NOLD_VEL  $MA_LOAD_TRQ  $MD_LOAD_TRQ  $MAX_TRQ_MGN  $MA_GRAV_MGN  $MA_STAL_MGN  $MA_BRK_MGN  $MA_NOLD_MGN  $MD_GRAV_MGN  $MD_STAL_MGN  $MD_BRK_MGN  $MD_NOLD_MGN  $PTH_GRV_MGN  $PTH_STL_MGN  $PTH_BRK_MGN  $PTH_NLD_MGN  $DYN_FRC_MGN  $MR_NOLD_TRQ  $R_ACC_MGN  $R_DEC_MGN  $R_LONG_MGN  $J_ACC  $J_DEC  $DT_MGN  $SP1  $SP2  $SP3  $SP4  $SP5  $SP6  $SP7  $SP8  6�TBJ_GRP_T   $$TBJ_ACCEL1   	$TBJ_ACCEL2   	$ASYM_PARAM   $TB_PARAM 2 	$SHORTMO_SCL  $LONGMO_SCL  $MIN_ACC_SHM  $MIN_ACC_UMA  $SHORTMO_MGN  $LONGMO_MGN  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2J_UPR_ANG  $J2J_LWR_ANG  $J2J_UPR_MGN  $J2J_LWR_MGN  $INERTIA_VIB   $INERTIA_VI2   $IV_UNIT  $IV_UNIT2  $R_F2JACC  $R_F2JDEC  $R_F2JLONG  $MIN_F2JACC  $MIN_F2JDEC  $MIN_F2JLONG  $MIN_ACRJ_S  $MIN_ACRJ_L  $MIN_PAYLOAD  $HVAL   $HMGN   $HAXS   $FLEX    ��TCPPIR_T    $ENABLE_TCPP  $TCDELAY   �|�TCPPSPEED_T  X $TCDELAY_MON  $VSPEED  $SPEED  $ACCEL  $TIMESTAMP  $PROG_SPEED  $MOTYPE  �TCPP_CFG_T 	 | $NUM_TCPPSEG  $GROUP_NUM  $TCPP_TIME  $WARNING_ENB  $OTF_TIM_ENB  $DEBUG_TASK  $DEBUG_MAIN  $TCPP_CMP_SW  ��TCPSPDCFG_T 
 � $TCDELAY  $HEARTBEAT  $SETUP_CFG  $SPD_MARGIN  $DEBUGFLG1  $DEBUGFLG2  $SPARE_STR1 $SPARE_STR2 $SPARE_LONG1  $SPARE_LONG2  $SPARE_REAL1  $SPARE_REAL2  }�TCPSPDOUT_T  p $ENABLE  $TARGET_TYPE  $TARGET_IDX  $MIN_VALUE  $MAX_VALUE  $MIN_SPEED  $MAX_SPEED  $GROUP_NO  �TP_THR_TABLE  $ $THR_ENB  $DI_NO  $DO_NO   #`�THR_CFG_T  0 $MAX_IO_SCAN  $MIN_SCAN_TI  $SCAN_TIME  ��TIMER_T  � $COMMENT $TIMER_VAL  $STR_EPT_IDX  $STR_LIN_NUM  $END_EPT_IDX  $END_LIN_NUM  $TID_NUM  $DUMMY13  $PS_OVERFLOW   $OVERFLOW  $FLAG_TYPE  $FLAG_IDX  $GLB_TMR_ENB  $GLB_TMR_STR  �TORQCTRL_T  X $DEBUG  $GRP_STT   $SBR_PAM21_V   T$SV_ERR_MOD   $SV_ERR_CLR   $ACTION  �TPGL_VIEW_T  4 $X  $Y  $Z  $WZ  $P  $R  $CAMERA   @�TPGL_UVIEW_T   $NAME $GIF }$VIEW ��TPGL_CAM_T  L $NAME $ID }$FID E$GIF }$NEARPLANE  $FARPLANE  $DISTANCE   ��JOG_RAD_T   $JOINTS   	��TPGL_MSET_T    $NAME E$ID }$TIMECONST  |�TPGL_CONF_T � $MOUNT ?� $LOCK_FOLLOW  $DBGLVL  $GLDBGLVL  $TEST_XML }$TEMPINT   $TEMPSTR ?� $USER_VIEWS 2 $CAMERAS 2 $TEMP_LOCS 2 $SCENE_VIEW 2  $KAREL_TMO  $TPDRAW_TMO  $JOG_VECLEN  $JOG_RADIUS 2 $CHECK_TOOLS  $CHECK_VIS  $REG_VIS32  $REG_VIS64  $MACHSET 2 $CONT_IDX  $DUMMY29  $VISIBLE   @$RAIL_BOXES   $ROBOT_XML ?� $SHOWWARN   $PS_CONTROLM   $CONTROLMAX  $CONTROLMASK   $FP_TO_FK ! ��TPGLMACH_T   $JOINTS   	X�RECLOC_T   $SLOTS !   ��TPGL_OUT_T  X $VIEWS 2 $SELECTED ?� $PIP_XML }$NODEVIS   @$MACHINES 2 $RECORDEDLOC 2 ��TPP_MON_T  D $GLOBAL_MT  $LOCAL_MT  $MON_NUM  $GMON_TID  $SYSMON_ADR  �TPSTRTCHK_T  , $ENABLE  $ALLOW_NAME $ALLOW_LINE   ��TPVWVAR_T  � $TPVIEW_ENB  $PREV_RTN  $EDIT_RTN  $VSHWRK  $DEBUG  $DISPLAY  $INDENT1  $INDENT2  $HEAD1 $HEAD2 $EDIT_KEY  $TCPSPD_KEY  $JMPCALL_ENB  `�TRACE_CFG_T  D $ENABLE  $ITEMS  $CHANNELS  $DEBUG  $TICKS  $MIN_MM  ��TRACE_CHNL_T  @ $ITEM_NUM  $TCP_GP_NUM  $VISIBLE  $STYLE  $COLOR   ��TRACE_ITEM_T  t 
$PRG_NAME %$VAR_NAME =$DESC !$UNITS $TYPE  $IO_TYPE  $PORT_NUM  $SQUARE  $SLOPE  $INTERCEPT  ��TSCFG_T  $GRP_MASK  $MODE_MASK  $STATUS  $OPT_VAL  $SIZE  $FNAME_TYPE  $PS_PROC   $PROC  $OUTPUT  $OUTPUT_DONE  $AXS_MSK_ENB  $AXIS_MASK   $CUR_RECTIME  $TOT_CHN_NUM  $MINFREQ_US  $SETFREQ_POW  $LPARAM   
$FPARAM   
$PATH_NAM $DUMMY19  $DUMMY20   P�TSR_GRP_T  l $MR_MAX_TRQ   	$MR_STAL_TRQ   	$MR_BRK_TRQ   	$MR_BRK_VEL   	$MR_NOLD_VEL   	$MA_LOAD_TRQ   	$MD_LOAD_TRQ   	$MA_GRAV_MGN   	$MA_STAL_MGN   	$MA_BRK_MGN   	$MD_GRAV_MGN   	$MD_STAL_MGN   	$MD_BRK_MGN   	$MJ_ACC_MGN   	$MC_ACC_MGN   	$MC_STAL_MGN   	$MC_BRK_MGN   	$MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	��TSSCB_T ! h $DSP_NO  $DSPAX_NO  $DATA_SEL  $OUT_CHANNEL  $ADDRESS  $BIT_SHIFT  $USE_2CH  $MONITOR  �TXSCREEN_T " $ $DESTINATION }$SCREEN_NAME  ��REQ_DATA_T # T $ERR_TYPE  $ERR_GRP  $ERR_AXIS  $AXIS_TYPE  $ERROR_DIST  $ERR_TIME   ��UECFG_T $ � 	$CHK_VERSION  $RSM_CHK_ENB  $UNEXCEP_ENB  $RSM_THRS_R  $RSM_THRS_L  $UNEX_THRS_R  $UNEX_THRS_L  $REQ_COUNT  $REQ_DATA 1# 
�UEGRP_T % 0 $ERR_COUNT  $PROGMTN_FLG  $CURR_POS   	��UI_MENHIS_T & 8 $HIST_HEAD  $HIST_ENTRY ?� $DUMMY2  $DUMMY3  \�UI_MOUSE_T ' @ $ACTION  $BUTTON  $ROW  $COLUMN  $TIME  $RESERVED  �UI_PANEDAT_T ( � $PAGEURL }$FRAME )$HELPURL }$PARAMETER1 )$PARAMETER2 )$PARAMETER3 )$PARAMETER4 )$PARAMETER5 )$PARAMETER6 )$PARAMETER7 )$PARAMETER8 )$INTERVAL  $PANESTATE  $DUMMY14  $MOUSE '�UI_USRVIEW_T ) < $MENU $CONFIG $FOCUS $PRIM m$DUAL m$TRIPLE m�UNDO_CFG_T *  $UNDO_ENB  $WARN_ENB  ��USER_INFO_T + 8 $USR_PROG %$TASK_ID  $USR_POSIDX  $USR_PR_USE  �USER_TOOL_T , 4 $X  $Y  $Z  $W  $P  $R  $TOOL_NUM  ��USER_UFRAM_T - 4 $X  $Y  $Z  $W  $P  $R  $UFRAME_NUM  �USER_OFFST_T . D $TOOL_OFST 1, $UFRAME_OFST 1- $GUN_WIDTH   $ENB_SUBNUM   
�USRTOL_GRP_T / @ $DIST_TOL  $ORNT_TOL  $RAUX_TOL  $TAUX_TOL  $ENABLE  �VCCM_CFG_T 0  $SC36MFB1ENB   !��VCMR_CAM_T 1h $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DETECT_TYPE  $DRIVE_TYPE  $SET_VTCP  $DEBUG_CODE  $DMY_UBYTE  $CAMERA_NAME %$DISTORTION1  $DISTORTION2  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $HANDEYE  $EXPOS_TIME  $NUM_MUL_EXP  $FOCAL_DIST  $GD_SPACING  $TRGT_DIST  $TRGT_W  $TRGT_P  $TRGT_R  $NUM_RETRY  $UTOOL   $�VCMR_TRGT_T 2  $TARGET_PNT   A<�VCMR_CRPR_T 3 d $AXIS_FLAG   	$NUM_AXS_REP  $SWING_ANG   $NUM_MS_POSE  $BASE_POSE   	$EVALUE_IDX   <�VCMR_CHKM_T 4 @ $EVALUE_IDX  $MAX_MS_ERR  $MEAN_MS_ERR  $WORST_POSE  ��VCMR_MRCV_T 5 � $ORG_MST_CT   	$ORG_UFRAME   $ORG_REF_POS   	$ORG_REF_CT   	$RCV_ANG_PAM   	$NEW_MST_CT   	$NEW_UFRAME   $NEW_REF_POS   	$NEW_REF_CT   	$EVALUE_IDX  $MAX_RC_ERR  $MEAN_RC_ERR  $WORST_POSE  $MASTER_TIME  $DEBUG_MODE   (�VCMR_GRP_T 6 � $STAT_FLAGS  $MENU_CODE  $GROUP_NUM  $UTOOL_NUM  $CAMERA 1$TARGET_ID 22 $CREATE_PRG 3$DATA_ID  $CHK_RESULT 4$RECOVERY 5$EXT_INT1  $EXT_INT2  $EXT_INT3  $EXT_INT4  $EXT_REAL1  $EXT_REAL2  $EXT_REAL3  $EXT_REAL4  �VISION_CFG_T 70 &$DATA_PATH  $DATA_CACHE  $LOG_PATH  $LOG_EXPATH  $LOG_TIMEOUT  $MC_LIMIT  $FR_LIMIT  $TD_LIMIT  $DEBUG_MODE  $HOST_NAME  $COMM_PORT  $ROBOT_NAME  $FLAGS  $MAX_PAGES  $MIN_VPOOL  $VPOOL_SZ32  $VPOOL_SZ64  $VPOOL_SZ128  $VPOOL_SZCAL  $VPOOL_LIM  $VPOOL_WAIT  $TMPPOOL_LIM  $FAILIMG_IDX  $LOADIMG_IDX  $NUM_IMREGS  $IMREG_SIZE  $GPM_CANDMAX  $NUM_ASYNBUF  $NUM_VRTDBUF  $VRTDBUF_SIZ  $TOLE_2D_Z  $TOLE_2D_WP  $PC_SETUP  $LOGQUE_MAX  $ECCU_RETRY  $VEMT_PATH  $VEMT_LIMIT  $VIRCIMG_SIZ  \�VISION_GRP_T 8  $BACKLASH   	�VLEXE_CFG_T 9 D $ENABLED  $DATE  $FLDR_INDEX  $FILE_INDEX  $REC_INDEX  x�CUSTOMMENU_T : $ $TITLE $PROG_NAME %$OPTION  �VSHIFT_CFG_T ;` $DATA_NAME 	$CAMERA_NAME %$EXPOSURE  $WIN_RADIUS  $WIN_POS_X  $WIN_POS_Y  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $LIM_DIST  $LIM_ANGLE  $LIM_TILT  $LIM_SCORE  $LIM_CNTRST  $WARN_DIST  $WARN_ANGLE  $WARN_TILT  $WARN_SCORE  $WARN_CNTRST  $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DUMMY23  $USED_CAMTYP   |�VSMO_CFG_T <  $ENABLE  $ADJUST_TIME  �WAIT_DATA_T =  $PROG_NAME %$LINE_NUM  �WV_AXSRST_T >   $AXIS_MASK  $THRESHOLD    ��ZABC_GRP_T ?  $ZABC_MODE   
 ��ZMPCF_GRP_T @   $ZMP_ENB  $ZMP_DMY_LNK   
h�ZMPOS_GRP_T A � $M_POS_ENB  $CMCMD_SCL  $CART_MCMD   	$P_ACT $J_ACT   	$P_DES $J_DES   	$P_DES2 $J_DES2   	$UXWPR_ENB  $UXEUL_ENB  $UXWPR_ACT   $UXWPR_DES   $UXEUL_ACT   $UXEUL_DES    ��ZP_CFG_T B  $ENABLE  $DEBUG  t�ZP_CYLINDER_ C 8 $RADIUS  $HEIGHT  $PROG_NAME ?( $LINE_NUM    ��ZP_GRP_T D � $OPTIONS   
$BREAK_TIME  $WORK_SHIFT  $ENABLE  $RV_LIFE   	$SHIFT_OVC   	$PART_ID  $OPTM_RATE   
$MAX_I_RATE  $MAX_DI_RATE  $TRACE_ENV  x�ZP_SPHERE_T E , $RADIUS  $PROG_NAME ?( $LINE_NUM   ��$TBC_GRP 2������� d � �?    	 HD)�?�  ?�  ??D�??D�?%�'?�  ?�  D)�B:ff                                D)�?�  ?�  ?333?333?��?�  ?�  D)�ByP                                D)�?�  ?�  ??D�??D�?%�'?�  ?�  D)�B�+�                                C?�  ?�  ?D�?D�?D�?�  ?�  CA��C&ff                                C?�  ?�  ?rw�?rw�?rw�?�  ?�  CA��C�I                                C?�  ?�  ?rw�?rw�?rw�?�  ?�  CA��C+�                                @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  ?�  ?�     �   �	V3.00     	rb21      	****      	�                              ?g!�?�     X   `?�  ?�                                            ?���Cz                                          ������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  �������������������������������������$TBJCFG �������                 �                                     �                                                 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                              	                                      	                                      	                                      	                                      	                                                                                      	                                      	                                      	                                         ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������                                             �$TBJOP_GRP 2�������  ?���C     	����������������������������$TBJ_GRP 2������� � 	 ����X�       	 �X^ �,X        @   ?�   	 �D)�D)�D)�C2
C랔        ?�  ?�  ??D�??D�?%�'?�  ??D�??D�?%�'?�  ?:p�?:p�? �U<p�SD)�>���?'!�?'!�B���B
�n    ?�                              D)�D)�D)�C2
C랔        ?�  ?�  ??D�??D�?%�'?�  ??D�??D�?%�'?�  ??D�??D�?%�'<?D)�?�?M�?M�C��B���    ?�                              D)�D)�D)�C2
C랔        ?�  ?�  ??D�??D�?%�'?�  ??D�??D�?%�'?�  ??D�??D�?%�';�ŗD)�>���?'!�?'!�C+�B�+�                                    CCCC���C�p�        ?�  ?�  ?s33?s33?s33?�  ?s33?s33?s33?�  ?D�?D�?D�;���CA�?@�??s�r?s�rCk�B���                                    CCCC���C�p�        ?�  ?�  ?rw�?rw�?fff?�  ?rw�?rw�?fff?�  ?rw�?rw�?rw�;�?)CA�?'!�?ZT�?ZT�C4+�B�$�                                    CCCC���C�p�        ?�  ?�  ?fff?fff?fff?�  ?fff?fff?fff?�  ?rw�?rw�?rw�;l�CA�?333?fff?ZT�CW�C+�                                    ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      C�         �   �?�  ?�  	V3.00     	rb21      	****      	�                                F�� F�. G
� G(� GG� Ggs G�� G�v G�^ G���G�@�G�; G쑀G�C�H	(�H� H��H&��H1�H;y�  F?� FM4 Fj0 F�` F�v F�V F� G> G7� GZj G�l G���G���G�� G�� G���HS@H��H0) HB�@=L��<�?�  ?�  ?�     @   X   `?�  ?�                                                          ?�  @   ?�  ?�                               	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  �������������������������������������$TCPPACTSW  ������    �$TCPPIR �������   CH  �$TCPPSPEED ������ CH                      U$�        �$TCPP_CFG 	�������                          �$TCP_SPD_CFG 
�������     dI   :�o        �              �                              �$TCP_SPD_NUM      ����   
�$TCP_SPD_OUT 2������� 
                                                                                                                                                                                                                                                                                                              �$TCZEROSPD              �$TESTPARS  ������   �    �$THRESTABLE 1�������                                                                                                 	           
                                                                      �$THRRDITABLE 1�������                                                                                          �$THRRDOTABLE 1�������                                                                                          �$THRSDITABLE 1�������                                                                                                                                                                                                                                                                                                                                                                                                   �$THRSITABLE 1�������                                                                                                             	           
                                                           �$THRTABLENUM  �������          �$THR_CFG �������   
   @   `�$TIMEBF_TTS         
�   �$TIMEBF_VER        
�   �$TIMER 1�������   8�                   �� ��  H��         �      �                   ͟� �  ��         �       �                     Y  ��         �       �                    g 	  ��         �       �                    <�� 	  ��         �       �                    $09 �  ��         �       �                   6�x���  H��         �      �                   :�x���  H��         �      �                   +�x���  H��         �      �                   W<	� ��  H��         �      �               B    x�x� ��         �       �                     �  �   ��         �       �               i     �  �   ��         �       �                     �  �   ��         �       �                n    �  �   ��         �       �               S_E    �  �   ��         �       �                      �  �   ��         �       �                      �  �   ��         �       �               �    �  �   ��         �       �               ST_    �  �   ��                   �               �9�    �  �   ��                   �               �    �  �   ��                   �               � �    �  �   ��                   �               �    �  �   ��                   �               u?�    �  �   ��                   �               _[_    �  �   ��                   �               '    �  �   ��                   �               ��    �  �   ��                   �               ��    �  �   ��                   �                ��    �  �   ��                   �               ��    �  �   ��                   �               w    �  �   ��                   �$TIMER_NUM        @�    �$TMI_CHAN          �    �$TMI_DBGLVL         �    �$TMI_ETHERAD ?�������  0000:e0:e4:13:cc:ae 0000:e0:e4:13:cc:af �                  0000:e0:e4:13:cc:b1 �$TMI_ROUTER !�������!ROUTER                            �$TMI_SNMASK ?�������  255.255.255.0     255.255.255.0     255.255.255.0     255.255.255.0     �$TOOLOFS_DIS         �    �$TORQCTRL ������                                       T                                                                                                                                                                                                                                                                                                                                                                                                                         �$TPE_DETAIL         �   �$TPGL_CONFIG ������  �?/cell/$CID$/grp1              ?�                                                                                                  �/cell/$CID$/grp2                                                                                                                  �/cell/$CID$/grp3                                                                                                                  �/cell/$CID$/grp4                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                             }�                                                                                                                                                                                  ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                    �User View 1           }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345 ���������������������User View 2           }�                                                                                                                              ���������������������User View 3           }�                                                                                                                              ���������������������User View 4           }�                                                                                                                              ���������������������User View 5           }�                                                                                                                              ���������������������User View 6           }�                                                                                                                              ���������������������User View 7           }�                                                                                                                              ���������������������User View 8           }�                                                                                                                              ��������������������� lCamera 1              }�                                                                                                                              E�                                                                      }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345             Camera 2              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 3              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 4              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 5              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 6              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 7              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 8              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 9              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 10             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 11             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 12             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 13             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 14             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 15             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 16             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   
   (  �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������                 �E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ����� @ ����������������������������������������������������������������  ��������  ��)frh:\tpgl\robots\r2000ix\r2000ib_210f.xml                                                                                                                                                                                                                 � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                            ���������     ����������������  88�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  �$TPGL_OUTPUT ������   ���?�              ?�              ?�                  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     }�                                                                                                                               @ ����������������������������������������������������������������  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  �  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8�����������������������������������������$TPOFF_LIM      ����   �$TPON_SVOFF         �    �$TPP_MON �������          2        �$TPSTRTCHK �������    �                  �$TPVTCOMPAT         �    �$TPVWVAR �������                   �                  �                       �$TP_DEFPROG %�������%FOLGE011                              �$TP_DISPLAY  �������    �$TP_INST_MSK  �������          �$TP_INUSER         �   �$TP_LCKUSER         �    �$TP_QUICKMEN         �    �$TP_SCREEN �������t_sc  �$TP_USERSCRN �������t_sc  �$TP_USESTAT         �    �$TRACE_CFG ������         	       
?�  �$TRACE_CHNL 2������ 	                 �                 �                 �                 �                 �                 �                 �                 �                 � �$TRACE_ITEM 2������  �%$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          �$TSCFG ������                 �  �                                                   
                                          
                                         UD1:\               ���$TSR_GRP 1 ������ � 	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678  �$TSSCB 2!������                                                                                                                                                                                                  �$TX_SCREEN 1"������ 
 �}ipnl/pnlgen.htm                                                                                                               Panel setup               }	index.STM                                                                                                                     
Robot Info e              }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          �$UALRM_MSG ?������� 
  �                              �                              �                              �                              �                              �                              �                              �                              �                              �                              �$UALRM_SEV  ������� 
   �$UECFG $������           @�  A�  A   B�     ! 
   �         @���X̌`  �          B���X̌`  �          B� X̌`  �         A� Ukys  �         A2�W�[|  �          B�ffX2+  �         B8�X�]  �          BɽfX�]  �          B� X�]  �         B	�X��$UEGRP 2%������  0       	 =���
�?
h=��뿽�/?�;�                    	 B�                                         	 B�                                          	                                     �$UI_DEFPROG ?%�������  (%MAKRO050 .......................0030  %MOTN005                               %�                                      %�                                      %�                                      %�                                      %�                                      %�                                      �$UI_INUSER  �������                                  �$UI_MENHIST 1&������  (   ��*/SOFTPART/GENLINK?current=editpage,UP023,1 ,4                                                                                     �-/SOFTPART/GENLINK?current=editpage,MAKRO050,1                                                                                     �'/SOFTPART/GENLINK?current=menupage,98,1 125,5                                                                                     �'/SOFTPART/GENLINK?current=menupage,71,1  1                                                                                        �-/SOFTPART/GENLINK?current=editpage,FOLGE125,5                                                                                     �'/SOFTPART/GENLINK?current=menupage,37,1 ,1 ,40                                                                                    �(/SOFTPART/GENLINK?current=menupage,381,1 11,33                                                                                    �-/SOFTPART/GENLINK?current=editpage,FOLGE011,5                                                                                     ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ���$UI_PANEDATA 1(������  	�}/frh/cgtp/doubdev1.stm 8981&action=100                                                                                        )prim                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ��    (�UD    }/karel/peeritp 1.stm m                                                                                                        )dual                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ��     �����}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}�                                                                                                                              )�                                          }�                                                                                                                              )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          ��������������$UI_POSTYPE  ������� 	                                    �$UI_QUICKMEN  �������                                  �$UI_RESTORE 1)������  ��                                             �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �$UI_SCREEN ?�������  u1sc  u2sc  u3sc  u4sc  u5sc  u6sc  u7sc  u8sc  �$UI_USERSCRN ?�������  u1ks  u2ks  u3ks  u4ks  u5ks  u6ks  u7ks  u8ks  �$UNDO_CFG *�������      �$UPDATE �������KS_24 �$USER_INFO 1+�������  0%FOLGE011                                    %                                               %                                               %                                               %                                               %                                               %                                               %                                               �$USER_OFFSET .�������                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                                   
                                        �$USEUFRAME         �   �$USRTOL_ABRT         �    �$USRTOL_ENB         �   �$USRTOL_GRP 1/�������  Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz     Cz  A�  A�  Cz     Cz  A�  A�  Cz     �$USRTOL_MENU            �    �$USRTOL_MSK         �    �$USRTOL_NAME %�������%�                                      �$VCCM_CFG 0�������    �$VCMR_GRP 26������               	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                    �$VISIONTMOUT        ��  ��$VISION_CFG 7�w`�x� FR:\VISION\DATA\                   �� MC:\VISION\LOG\                    UD1:\VISION\EXLOG\                  ' B@ �� ��     �                                                                                  �  =	 1- n6  -��         B@         ,             =���=���            MC:\VISION\TRAIN\                       �$VISION_GRP 28������  ( 	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���            �$VLEXE_CFG 9������    1-e            �$VMPHASE  ������          �$VSHIFTMENU 1:������ 
 <�              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���	LIVE/SNAP     %vsflive                               ���VISION SETUP  %vsfmenu                               ����              %�                                      ����$VSHIFT_CFG ;�������	�          %�                                        �5   @   �  @����       A�  B8  B  B�  Ap  Ap  B  A�  B�  B    �  ���������$VSHIFT_MEP        ���   �$VSMO_CFG <������    �z  �$WAITDINEND        �   �    �$WAITDINOK            �    �$WAITDINOUT        �   �    �$WAITDINST        �   �    �$WAITDINTIM       ��   �    �$WAITGINEND        �   �    �$WAITGINOK            �    �$WAITGINOUT        �   �    �$WAITGINST        �   �    �$WAITGINTIM       ��   �    �$WAITRELEASE         �    �$WAITTMOUT        ��  ��$WAIT_ACTIVE         �   �$WAIT_DATA =�������%$FOLGE011........................0006     �$WAIT_RDISP         �    �$WV_AXSRST 2>�������                                  �$WV_GRP_IR  ������ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �$ZABC_GRP 1?������  , 
        2                                 
        2                                 
        2                                 
        2                                �$ZMPCF_G 1@�������  0     
                                              
                                              
                                              
                                         �$ZMP_GRP 1A������  �      � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��  �$ZPCFG B�������        �$ZP_CYLINDER 2C�������  �          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZP_GRP 2D�������  � 
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�  �$ZP_SPHERE 2E�������  �      ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZZZ         ��    