��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�MC_CFG_T�   � $�'NUM_MSK�  $EXE�_TYPECME�M_OPTPN_�CNFCIF_C�Y:gSCN_T�IME E RESET_P�Do �LJ �HECK_�DSBLC $D�RA> ARGIN�CSTORJ �0&DEV. �d 	7OC'H�AR�ADD�S�IZORACBS�LO[ODKIO>KOCCPYC&|l /  L ���h99IDX���&L. � 
�EQPLH�RAT�TRKB�UF| ��UN_STATUS�sCU��MAX(�I����SNP_�PA�  �{ � ANNE��� OW CTION�_�PU�  � $BAUD��NOISYmNV�T1�#2�#3�$7_PR�T4P' �DATA�CQUwEUE� PTH[$�MM_��%&!RE�TRIESCAU�TO!R[��B�G � �ISP_�INFd�' CL�IMI� B5AD_ H C3H��#d6�#d6 �#d6�#W1� �#�4�#�4�#�4�" ��$$CLASS ? ����1��m���iFG0 ��5��� C�2��>!>!d��C\�3�  2�7	@d $DZO��WO�O {O�O�O�O�O�O�O_ _@_/_d_S_�_w_�_ �_�_�_�_�_oo<o +o`oOo�oso�o�o�o �o�o�o8'\ K�o����� ���4�#�X�G�|� k�����ď���׏� ��0��T�C�x�g��� �������ӟ���,� �P�?�t�c������� ���ϯ��(��L� ;�p�_���������ܿ ˿ ��$��H�7�l� [ϐ�ϴϣ������� �� ��D�3�h�Wߌ� {߰ߟ���������� �@�/�d�S��w�� �����������<� +�`�O���s������� ������8'\ K�o����� ��4#XG| k������/��0//4,�3IF �2CKP DX�D�G�%�@�@!�,�$"A�)�$�,��$�+JA@<(�!�()DY�(1�%/0�&I"<<�%<<�%<<�%	<;6E�55S1
'5F�(�(�1�!�!Q�;�"�!�<�� UH@��8G�(,L��5,K
F\L#E�"�8K�4k10'k5�@S��4�A��4R�3[�3*��4D�3C�@C�F7@C"H@DA�7�F�1U&_!_3_ E_n_i_{_�_�_�_�_ �_�_�_ooFoAoSo eo�o�o�o�o�o�o�o �o+=fas �������� �>�9�K�]������� ��Ώɏۏ���#� 5�^�Y�k�}��������şS/e"TYPE �2o+ (�3:�!d�6�|蟮1�ڞ�0L���ZA t����!��կ���b!�SNP_PARAOM o+ΥϯƧ�A'� S�̦�0[A �"�1l��1�!U&��) 4�