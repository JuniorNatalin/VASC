A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DRYRUN_T   � $DRYRUN_ENB  $NUM_PORT  $NUM_SUB  $STATE  $TCOL_SYSPT  $PMC_SYSPT  $GRP_MASK  $STEP_MOTION  $LOG_INFO  $TCOL_SAVE  $FLTR_EMPTY  $PROD_START  $ESTOP_DSBL  $POW_RECOV  $OPR_DSBL  $SAW_PROG %$INIT_PROG %$RESUME_TYPE  ��DRYRUN_PORT_  4 $TYPE  $FST_IDX  $LST_IDX  $STATIC_PORT  ��MIX_BG_T  4 $PROG_NAME %$MODE  $STATUS  $MODIFY_TIME  h�MIX_MKR_T   $LINE   $LINE_SIZE  `�MIX_LOGIC_T , $USE_FLG  $USE_MKR  $USE_TCOL  $USE_TCOLSIM  $NUM_FLG  $NUM_MKR  $NUM_BG  $NUM_SCAN  $MAXNUM_SCAN  $MINNUM_SCAN  $ITEM_COUNT  $PROC_TIME  $MAX_TMR_VAL  $TCOL_LINE $TCOL_ENB  $TCOL_SIM  $TCOL_STAT  $SAVE_IDX  $SAVE_LINE $TCOL_WARN  $BG_HITEM  $INST_CHK  �$$CLASS  ������   5    5�$DRYRUN  ������5�      c                        ����                   %VAGSAW                                %VAGTPINI                                 �$DRYRUN_PORT 2������5� c    "      $             d                   )     �                                             	  	                    �  �         �  �         �  �         �  �         �  �                    !  8         c  c         h  i         l  l         y  �         �  �         �  �         �  �                      	                      2         9  ;         A  P         a  x         �  �         �  �         �  �         �  �         �  �         �  �         �  �         �  �           !         )  +         C  C         H  I         L  L         Q  q         y  {         �  �         �  �         �  �         �  �         �  �         �  �         �  �         	  	         !  3         7  7         I  I         a  s         w  w         �  �         �  �         �  �                                 1  A         V  a         v  �       )   D   G       )   M   P       )   y   z       )             )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )           )  !  !       )  2  2       )  J  J       )  A  A       )  P  P       )  `  c       )  e  e       )  u  x       )  z  z       )  �  �       )  
  9       )  �  �       )  �  �                                                                                                    �$DRYRUN_SUB ?������5�  FOLGE         UP         0  MAKRO         SUCHL         BIN1        D�$MIX_BG 2������5�  4%MAKROSP1                                    J�]P%MAKROSP2                           </t      J�]Q%MAKROSP3                           h=3      ����%MAKROSP4                           5-1      ����%MAKROSP5                           ="4      ����%MAKROSP6                                    ����%MAKROSP7                           ame      H��%MAKROSP8                            �      J�]Q�$MIX_LOGIC ������5�                  �              X  ����  s2tq* q* q* !q* _q* `tq* q* !q* _q* `t                                                                                                                                                                                                                         ����  s2tq* q* q* !q* _q* `tq* q* !q* _q* `t \ttq�tt�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������             �$MIX_MKR 2������5 �  * dss
Mtr
 t
 t                                                                                                                                                                                                                                              * dsu
Mqu
Ot                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       * ds
 +q
 -t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             * ds
 q
 q
t                                                                                                                                                                                                                                                * ds
Cqu
Dq
Equ
Fq
Gqu
Hq
Iqu
Jt                                                                                                                                                                                                                 2  *  dsu
Cq
Dqu
Eq
Fqu
Gq
Hqu
Iq
Jt                                                                                                                                                                                                                 2  * !dsu
Kq
Lt                                                                                                                                                                                                                                                    * "ds
Kqu
Lt                                                                                                                                                                                                                                                    * #ds2 t                                                                                                                                                                                                                                                          	  * $ds2 t                                                                                                                                                                                                                                                          	  * %ds2 t                                                                                                                                                                                                                                                          	  * &ds2 t                                                                                                                                                                                                                                                          	  * 'ds2 t                                                                                                                                                                                                                                                          	  * (ds2 t                                                                                                                                                                                                                                                          	  * )ds2 t                                                                                                                                                                                                                                                          	  * *ds2 t                                                                                                                                                                                                                                                          	  * +ds2 t                                                                                                                                                                                                                                                          	  * ,ds2 t                                                                                                                                                                                                                                                          	  * -ds2 t                                                                                                                                                                                                                                                          	  * .ds2 t                                                                                                                                                                                                                                                          	  * /ds2 t                                                                                                                                                                                                                                                          	  * 0ds2 t                                                                                                                                                                                                                                                          	  * 1ds2 t                                                                                                                                                                                                                                                          	  * 2ds2 t                                                                                                                                                                                                                                                          	  * 3ds2 t                                                                                                                                                                                                                                                          	  * 4ds2 t                                                                                                                                                                                                                                                          	  * 5ds2 t                                                                                                                                                                                                                                                          	  * 6ds2 t                                                                                                                                                                                                                                                          	  * 7ds2 t                                                                                                                                                                                                                                                          	  * 8ds2 t                                                                                                                                                                                                                                                          	  * 9ds2 t                                                                                                                                                                                                                                                          	  * :ds2 t                                                                                                                                                                                                                                                          	  * ;ds2 t                                                                                                                                                                                                                                                          	  * <ds2 t                                                                                                                                                                                                                                                          	  * =ds2 t                                                                                                                                                                                                                                                          	  * >ds2 t                                                                                                                                                                                                                                                          	  * ?ds2 t                                                                                                                                                                                                                                                          	  * @ds2 t                                                                                                                                                                                                                                                          	  * Ads2 t                                                                                                                                                                                                                                                          	  * Bds2 t                                                                                                                                                                                                                                                          	  * Cds2 t                                                                                                                                                                                                                                                          	  * Dds2 t                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              * _ds
�qu
�q
�q
�qssu
�q
�tr�tqu
qu
q�t                                                                                                                                                                                                   @  * `ds2tJqu
Lqu
Kq
Mqu�qs)Arskq) �trsq) �ttt                                                                                                                                                                                                  	  * adss
�q�r)8tq
BqBqu) Hqu) Iqs) Zr) \tt                                                                                                                                                                                                          9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          