��   ɋ�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_CPC_�T   � �$COMMENT� $ENA�BLE  $�MODJGRP_�NUMKL\ � $UFRM�\] _VTX �M �   $Y��Z1K $Z2��STOP_TY}PKDSBIO��IDXKENBL?_CALMD�&}S. � 8�J\TC�u
SPD_LI_����COL�&Y0 � � !CHG�_SIZ$A�P7ECDIS � � �7�C�����Jp 	�J �� ��"��$�'"_SEs��xSTAT/� D $FP_�BASE �$LINK`$!��j&_Vs.Hs# �(&J- ���ZAXS\UPR:LW�'CU�� `�$� | 
�/�/�/4�??j&ELE�M/ T $1Uc c1j"NO�7�0�a3UTOOi�2H�A�4�� $DA{TA" &e0   @P:�0� 2 
&PNP% ��P!U*.n   oFSyCjHrB� zB(�F�D(�1�R5C�DROBOT��H�CQBo�E�F$CUR_"�B��SETU�	 l|� �P_MGN�INP_ASS�  @�� �3�8"7GP@ U�>VhSP!�T&T1�
@B\8�8�T= 0 P�+ Kec1VRFY�8�T$5&1�� ��W��1k$R�0TPH/ ([ �#A�#At�#A3tBOX/ 8�0����Г`bo%ch�TUI}R�0  ,[ ��62`ERa02 {$k` �a�_S�b�fZN>/ 0 [9&02� arZ_� ��_� tu0  @��A�Yv	�on \��$$CL,P  O����q��Q��wQ�$' 2 �u�Q   ���q���b0�p�}�p��~� 4�F���m����� �ǏُL������� E���i�{���$� 6��Z�����A��� Ɵ؟��������2�� V�h�z�+���O�a�ԯ ����
�@�Ϳ���� v�'Ϛ����п^ϓ� �����<�N���r�� 5�Gߺ�k����ϡ�� ������\��ߒ�C� ��g�y��ߊ��"�4� ��X�	����?����� ��������0���T� f�x�)��M_��� ���>�t %���m\�� �:L�p�3/ E/�i/��q//�/ �/�/Z/?~/�/A?�/ e?w?�?�/�? ?2?�? V?OO�?*OOO�?�? �O�?�O�O.O�OROdO vO'_�OK_]_�O�_�O __�_<_�_�_r_#o �_�_�_ko�_�o�oo �o8oJo�o�o1C �og�o�o"�� �X	�|���O� u�������0��T� ��)���M���ҏ�� ������,�ʟ�b�t� %���I�[�Ο��� �ǯ:����p�!��������i�ܯ�������$DCSS_CS�C 2I�ɱ�Q  D ���@���&���J� \�n�=ϒϤ϶υ��� ������"�4��X�j� |�Kߠ߲��ߓ����� ���0�B��f�x�� Y����������� ��>�P�b�1�����g������������GR�P 2ɻ ��	��cN�r ������ ;&Kq\��� ���/�%//I/ 4/m/X/j/�/�/�/�/ �/�/?�/3??W?B? {?f?�?�?�?�?�?�? �?OOAO,OeOPO�O �O�O|O�O�O�O�O_ __O_:_s_�_T_f_ �_�_�_�_o�_'oo 7o]ooo>o�o~o�o�o �o�o�o�o5
STAT 2ɹ�Y�,8�?��k?&L�?�I?Q���NW��%�=��K?���RhC�|IC�t�D�N:ɱ�,p8xr52?5����nW4nW�?�  �q���p4��ZC\?�UC\���ɱ^xq�����p;�p�=�  ^�p��5��yÞp̾�RD>	@�v����(�0?D�����p/�
nr�
�@�,�$����ђ�L�Z�Di S�v=�"��+@�?8G��@��@�)H��?Q����pv�p�C��Ą��D�h���u|p��p�p?��y�?Ns>�%�ѽ�o���?Ri��z� �́ɵ��ɵ�J� \�:������z�p��� ���ş�ٟ�%�� !�3�E�W�y�{����� ٯ�v���d��H�Z� 8�~�����䯺���ƿ �ڿ��&��2�\�F� hϒ�|ώ��ϲ�p�
� ���@�R�0�v߈�f��Ѐ�?&M�?��x����q���&[=��?����R[C��~kC�w2D�M��{�p/r�p�j�p=�s����s���p�{���p�p��pw�p�z�6��Þo�@���� ���T���?D��p#�߾<��
�l�+�$�G�ёK����Di!	X�����+?�?8HU�l�l�(t�Fx�����~��UC�U|��ǌ�1����֟����਀{>��&^���5���?R\�� �߸���l�>�P�.�t� ��d������������� ��(R<N� r������� 6H��l~\�� ����/�/ 2/4/F/h/�/|/�/�/ �/�/�/$.?@?�d? v?T?�?�?�?����� ������&�8�J�\� n����������O �?�?"��?n_�?^_�_ �_�_�_�_�?o�/ "oLo6oXo�olo�o�o �o�o�o�o�o$�_ fxV����� �_8��D�.�P� z�d�v�������ΏЏ ��.��^�p���� ����ʟܟ�?,_>_�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ��R_��������Կ ���
���<�F�� R�|�fψϲϜϾ��� ������*�T�>�� ��迆����߼��� .�h�>�D�J�t�^�� ����������� � �L�6��ߎ���~��� ��������\�n�,� >�P�b�t��������� ί����(�:�$ 6H�������/ �(/:/ �J�d/n�`/ �/�/�/�/�/�/�/? ?$?N?8?Z?�?v��? �?/�?�?�?O2OL/ ^/�?nOt?zO�O�O�O �O�O�O_�O_F_0_ R_|_f_DO�_O�_�_ o�_*o<oz��\ n������� �"lFXjTo foxoo���"�4� �X�j�PO�_���_�� ʏ��Ə ����� � 2�T�~�h������_� ��H��,�
�P�b�|� ����ʟ��������� 
����@�*�L�v�`� ����ҟܿ�@���$� �4�Z�8Ϫ���o �o�o�o�o�o�o
 .@R�v��߄� ���J��.��R�d� B������� �����0��<�f�P� b�����������z� &J\:���� ���������( $FHZ|�� ��//pB/T/ 2/x/�/t����ߪϼ� ��������(�:�L� ^�p߂ߔߦ߸��ߴ/ �/ �/LO�/\O�O`O rO�O�O���O� _ *__6_`_J_l_�_�_ �_�_�_�_o�_�ODo Vo4ozo�ojo�o�o�O o�o�_�o".X Bd�x���� ���o<�N�,�r����b������e�$DC�SS_JPC 2��eQ G( D��%�� $�6�H��l�~���_� ��Ɵ�������ݟ2� D�V�%�z�����m�¯ ԯ毵�
�����R� d�3�������{�п� ��ÿ�*����`�r� AϖϨϺω������ ��&�8�J��n߀�O� a߶��ߗ�������� 4�F�X�'�|��]�o� �����������B� T�f�5�������}��� ������,��Pb tC������ ��(:	^p� Q����� // �6/H//)/~/�/_/ �/�/�/�/�/? ?�/@D?V?%?7?#�؅S���@BS �HALT�?u5u? � )�=����?�?�4�?�?O�6! O2ODO�6`OrO��O�6�A�O�O�O�3�O�OC_�6 _2_�_B�6`_r_�_�6	�_�P��_ox?$��_Eo o*o{oNo�oro�o�o �o�o�o�o�oA& wJ\n���� ���=��a�4��� X�j�����ɏ���֏ �9���0���T�f� ����������ҟ�"� G��,�}�P���t�ů ������ί	��C�� (�y�L�^�p������� ��ʿܿ�?��$�b� ��Z�lϽϐ��ϴ�� ����;��I�2߃�V���?_MODEL ;2�;xt�i�W
 <m�c�:�H�J"����X�/�A� S�e�w������� ������+�=���a� s��������������� g�P��+�o� �������L #5�Yk}�� � /��6///1/ C/U/g/=�/a�/�/ ?�/�/D??-???�? c?u?�?�?�?�?�?�? �?@OO)OvOMO_O�O �O�O�O�O�O�O�/�/ �/__�_�Om__�_ �_�_o�_�_8oo!o 3oEoWoio�o�o�o�o �o�o�o�ojA S�;_M_{��u ����+�x�O�a� ����������͏ߏ,� ��b�9�K�]�o��� ������ɟ���� �p��Y�k������� �ůׯ$�����l� C�U���y���ؿ���� ӿ ���	�V�-�?ό� '�9�K�yϋ�a����� .���d�;�M�_�q� �ߕ��߹������� �%�7�I��m���� ������&������ ��E�W���{������� ��������X/A �ew���� ��B+=�� 7�ew���/� /P/'/9/K/�/o/�/ �/�/�/?�/�/�/L? #?5?�?Y?k?�?�?�? �?�O��?�?ZO1O CO�OgOyO�O�O�O�O _�O�OD__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o�?�o#OQo co�o�o�o�o�o %7�[m�� �����8��!� n�E�W�i�{�����uo ���oǏُF��/�|� S�e�w�ğ������џ �0���+�x�O�a� ������䯻�ͯ߯,� ������=�O��� 7�����ɿۿ�:�� #�p�G�Y�k�}Ϗϡ� ������$�����1� C�Uߢ�yߋ���s��� ����2���-�?�Q� c����������� ����d�;�M���q� ������������ N����);�#� ����&�\ 3EW�{��� �/��/X///A/ �/e/w/�/_q��/ �/�/??f?=?O?�? s?�?�?�?�?�?O�? OPO'O9OKO]OoO�O �O�O�O_�O�O�O�$��$DCSS_P�STAT ����cQQ?    t_�Z r_ (�_�_�WpkPkP�_�_ l cdP��P;_4oFo�)"ocUcUdovo�TTSETUP �	cYB�&T�#��!�dOYT1SC �2
�j`�!Cz��#/}�eCP [R�l�� DSo z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ��.h%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛ���������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� ����}����������� ����1CUg y������� 	-?Qcu��������Z�D �/*/</�/`/r/�/S/ �/�/�/�/�/??�/ 8?J??[?�?�?a?�? �?�?�?�?O"O�?FO XOjO9O�O�O/}O�O �OoO__0_�OT_f_ x_G_�_�_�_�_�_�_ �_o,o>ooboto�o Uo�o�o�o�o�o �o:L�O)�� ���� ��$�� H�Z�l�;�����q��� ؏ꏹ�� �2��V� h�z�I�������� ��_՟.�@�ǟd�v� ��W�����Я����� ��<�N��_����� e���̿޿����&� ��J�\�n�=ϒϤ�s���$DCSS_T�CPMAP  �������Q @ ~�J~�~�~���~�U~�~�~�	g�W  ~�~�~�U~�~�~�~�U~�~�~�~��~�~�~�~��~�~�~�~��~�~� ~�!~�"�~�#~�$~�%~�&�~�'~�(~�)~�*�~�+~�,~�-~�.�~�/~�0~�1~�2�~�3~�4~�5~�6�~�7~�8~�9~�:�~�;~�<~�=~�>�~�?~�@��UIR�O 2�����$��"�4�F�X� j�|��������������0�B�T�}� �}����������� ��1CUgy �����^���� �-?Qcu�� �����//)/ ;/M/_/��/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�?��?v/O��UIZNw 2��	 �����PObOtOy�KO�O �O�O�O�O�O_�O0_ B_T__x_�_�_k_�_ �_�_�_�_o,o�_Po boto�oIo�o�o�o�o �o�o:L^- ���i���� �$�6��Z�l�~�M� ����Ə؏�����ݏ�2�D�V�O��UFRwM R���� �џ���ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߒ��߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s��ߗ��� ��������'9 K]o����� ���#5GYk���x��� ���//�B/T/ //x/�/e/�/�/�/�/ �/�/?,??P?b?y ��?�?I?�?�?�?O O�?:OLO'OpO�O]O �O�O�O�O�O�O�O$_ 6__Z_l_�?�_�_A_ �_�_�_�_o�_2oDo ohozoUo�o�o�o�o �o�o�o.	Rd {_��9���� ���<�N�)�r��� _�������ޏ��ˏ� &��J�\�sw