��   �A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG �DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��H�DwNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !���* D� $PRIMA�R_IG !$ALTERN1�<WAIT_TI|A ���FT�� @� LOG�_8	�CMO>�$DNLD_FI�:�SUBDIR�CAP� D���8 . 4� H��ADDRTY�P�H NGTH�����z +L�S�&$RO�BOT2PEER�2� MASK4M�RU~OMGDEyV�� �RCM?�  $Z ��QSIZ�X��� TATUSWMAILSERV� $PLAN� �<$LIN<$�CLU���<$T�O�P$CC�&F�R�&�JEC�!��%ENB � A�LARl!B�TP��3�V8 S���$VAR9M O�N
6��
6APPL�
6PA� 5B 	7P�OR��#_�!�"A�LERT�&�2UR�L }�3AT�TAC��0ERR�_THRO�3US0�9z!�800CH- Y��4MAX?��R�DM*� $D�IS� ��S�MB�	"�BCA�$WI2�AIN4EXPSܣ!�PAR�
��0BCL�
 <�(C�0�SPTM3OU�4� WR�_H�uF �0@oC l5��!�"%�7,X�ECC�%� �VR�0UP� _D�LV�vE��S)No3 �O�B�X_S@~#Z_INsDE
B�QOFF� �~UR�YD���KT�   ts �!&PMON�r�SD��RHOU�#END�X�Q�V�Q�V�LOCA� Y$�N�0H_HE���TCPI"/ >3 $ARPz&�1F�W_\ �I!YF�P;FA~Lk0�1#�HO_� IN�FO7cEL	% �P K  !k0W�O�@ $ACCE� LV�K�2�H#ICE��` � ��$�c# ����q��
��
��$'0 u
U���F����It�Du�$� 2,{�a��r|}]p�� ,}��!q����r%r,z���0��AtDq�s`_  ,{�Krr����� ����̏ޏ����&��8��t� _FLTRs  v4s ���������{nx�,}2�{ZbSHw@D� 1,y  P��Atџ��� 2���V��z�=���a� ��ԯ�������߯@� �d�'�9���]����� ⿥��ɿۿ<���`� #τ�GϨ�kϡ����� ���&���J��V�1� ߤ�g��ߋ��߯�� ��4���	�j�-��Q� ��u��������0� ��T��x�;�q�������������wz _LI�� 1]�x!1E.10����01A>��255.y8&���Iu/26H@� \n���3��H%���
�4 &H�L^p��5�H �����6/H� </N/`/�r/L�RCj`�p�p!Pp%�ː�v� 'Q� ���.<(?]? o?B?�?�?�?�?�?�?��P�?O/OAO OeO wO�O�OZO�O�O�O�.�O��Lu-_\_�O�r_�_�_�_��}i�RConnect�: irc�T//?alerts�_�_ oo%o�Ul_QocouoЇo�o�o���� � �"<��d� DM�%s�~�$SMB 	���@o�/�C�v�`_CLNTw 2
�� 4#T-�\���� ���3��$�i�H� ����~�ÏՏ����N-M���n%�L�T��:�{��j������ǟ\�aN�1��m%172.+20� 4�3ӟ(v}������8����#�USTOM' �m3���0� ���$TCPIP�b�mX5 �TEL�e1�>2�H!TP!�#{�rj3_tp�dן # ��!KCL�諻���)u?!CRTB�0����2�!CO�NS�����smon���