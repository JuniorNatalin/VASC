��   v��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<�$1_8k����FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\9 ^75z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D��VCAX_�w A.  @ 5vFX0OR�@E ?NUM_SE238�_TO0Q�#RE_:� 2cT �+V>1 , $� �ME�vUPgDAT�wAXy_2 	�+VS5Q' 8<P��PnP;0k L\�R�PA�kQ�Q��+VM5Q  �$ISRTd 5+VG5Q { v��R2 
v�S2�T kR9�P 	��$U1SS  O����a����w�$' 1 �e� } �� 	 ����o�o�o�fZ�	�< �Fi���4 ��4R��o�oA,eP���xu}�a��}��l��s���ʀ��t��Jէ� �n�|�+�=�d�a��s� ���vB z����  B�����|� ����������K��_������.���o\��������pU0pgpx��d��1�C�U���=L���`���?�����@� ��͟ߟ���'�9��K�]�o������� ��e��̧��쯄d  2 ��/�A�S�e�w� ����������<�� ����1�C�U�g�y� �ϝϯ����`�a�o�� ����*�<�#�`�K� ��oߨߓ�y��ߡ�� ��&�q�5�G�n�k�}� �������������"� ��P�b�t������� ��������(: ��^p������ Eϯ��6HZ l~�����˿ �/ /2/D/V/h/z/ �/�/�/�/�/���/� �/.??R?9?v?a?�? �?�?�?���?�?OO <O'O�?]OoO�O�O�O �O3O�O�O_�O_J_ =�k_}_�_�_�_�_�_ �_�_oo1oCoUo |o�o�o�o�o�o�go io�o-#Tfx� �������� ,�>�P�b�t������� ��Ώ����/�(�� L�7�p�W������ʟ ����?�՟6�!�Z� l��O{�������ïկ Q����2�D�/�h�[_ ��������ѿ���� �+�=�O�a�s�5�� �Ͼ�������G���'� K�Ar߄ߖߨߺ� ���������m�J� \�n�����������������$FM�S_GRP 1�^� �>�H*~�G��G��H����H�'�I�}�J�ND��O�$�O]�+�K}�sKp���Iό�J�B� � ����~�A�������C�W�yA���C�SN�J���� �O���QB��P� L��/�L�$K�M���A7��?�����H*��G���G�NH����H�(�I}=�+�W
���������*� .� �$ 	RW�9�RkwRr��@R��Sy�@@U�I0VW�BċNkU�N�oEOmo$P�֬�P�KdQ�'�Q(;�Q�(^�Q(r�Q��JR) -R�-7iY�-Y�	��
�-��&�8 ����^9�a� ���RE�� ��D� �\vF�P��D���YFF�F���۷��G�с��*d�RE�h��P���2�7�ai�cͬa���j�?'���'8�2�>�(a���a�b>���?	�b���a��b���c0�a���@I�a�C�cg�"1s� �1�= 2�x�1_ ����0��0�4 ��
	 2�1 �2�� �A� ���7 2c �2�m 2p �2M 2�; W��ק rk �7����2���\s���U�V����
�U:���������UF�U]v������*����� A��{V.�����kv"�d��Z���Z�~N� i������� ik0�Z��w�Z�! i�Wu i�T�Z���Zļ�Z��%�[x�Z�� i�8�Z����Z�,7������7����������w������������w��������w�W�w΅�0���������0���}��w,�����ѻ}��?�?�?��?}��2'�  �M_�f�'�  ��  �  %_L  �_��_���  �4�D�����_��;@� W _��'@xKC�'p�4�  ��� ����������nG@&�_��_���;������_�����ύ  �_���A
�C47��k��'@���,�@�h���"@ e04�4��@��4�_B  �4� G@U�@�4��@�4��s@L�3�@�5�_�}@3�m�~��@k@m_Ф_�Ŭ4�P%@_Є�  �,�_Ћ�4�_Ж0@��D�ʔ@��@�w@2@@��@&P�e�o�@��_К@	K4������^���0@�����B@���
Qi�g��O�C-Q4�V�@ _��_��4�i�_�n@ �P K�@�>Av4��4�4�f�s@�4�r@��4��@ų4vPoo)o;oA`�3Yo�gco�o���B �@�b�aZ4� �d�a�e�a�i�i�g8��!�;��p���b-�$5����M&�>{O�p���`ɿ��W̿�f3���R��[��˿^>��XFp��3p��_N���1/p�#pb"?�X�>u��>t��^?�q>���?�^?��>��>t�NW>u>�>���>w>t��8>tU`>t�I�>tP�>t��x>#~>t��J>uI7��<�a�O�(��O�@�Hyc���񚾤�Z����l�����Oj^�O�0�p����i�O����Ol��Oh���pܿO�a�����O����O��7@��c�@�.:@�4�@�J@q��@��r�k@q�	@�7�@��2W@qc@q�e@�5`�گ@�8)3����@q@�+�D��Or���8���7��?�|��>�!?��?��>�����7�F�7��>��>�� ��7�N�7��7�7o��7���>��B�7��ѿ7�OrT����j'���d?R��@k��E?<�����@l���H�����@k��@l�ݾ�IE��������������<�@k���E8���#�	,($UP00	1�o� ��4��X� ?�Q���u�������� ϟ���B�)�f�M� �����������˯ݯ ��>�%�7�t�[��� ���ο���ٿ�(� �L��p�[ϔ�ϑ� �ϵ��������6�!� F�l�Wߐ�wߴߟ���������:�j Y�k�}���߳���T� �������1�C�U�g� &��������������� 	��-?Qc"� ���|��� );M_��� �x��/�%/7/ I/[///�/�/�/t/ �/�/�/�/!?3?E?W? ?{?�?�?.ʧBp?�? �?�?d?O/OAOSOO wO�O�O�OlO�O�O�O �O_+_=_O__s_�_ �_�_h_�_�_�_�[���1234567890o'e5�oIo9o mo]oyo�o�o�o�o�o �o�o!-5G{ k������� ���S�C�_�g�y� ��������ӏ���� �7�a���ﲟ�� �ӟ���0��T� ?�x�c�u�����ү�� ����,�#�P��_t� ������	����o�� �(��L�^�pς�A� �ϸ����ϛ� ��$� ��H�Z�l�~�=ߢߴ� ���ߗ���� ���D� V�h�z�9������� ����
����@�R�d� v�5������������� ��<N`r1 ����?�� 8J\n-�� �����/�4/ F/X/j/)/�/�/�/�/ �/�/�/?oc�9?Q� ]?M?i?q?�?�?�?�? �?�?OOO%O7OkO [OwOO�O�O�O�O�O �O�O_C_3_O_W_i_ �_�_�_�_�_�_�_o o'oQoAouou�?�o �o�o�o�o�o D /Aze���� �����@�7�d� v��/������Џ/�� ���*�<�N��r��� ��U���̟ޟ🯟� &�8�J�	�n�����Q� ��ȯگ쯫��"�4� F��j�|���M���Ŀ ֿ迧���0�B�� f�xϊ�IϚ������� ����,�>���b�t� ��Eߖ߼������� �(�:��^�p��A� �������� ��$� 6���Z�l�~�=����� �������� 2)? MeoYas��� ���'[ Kgo����� ���3/#/?/G/Y/ �/}/�/�/�/�/�/�/ �/?A?1?e?U?q?y?��1�$PLCL_GRP 1����1� �D�0�?� � �:]��?qg�9�O�:O%O^O IO�OmOO�O�O�O�O  _�O�>2_�OY_�O}_ h_�_�_�_�_�_�_�_ o
oCo*o$_vo8o�o 4o�o�o�o�o	 ?*cN�nho� |�x��)��M� _�J���n�����ˏ=��$VCAX_R�EF�0 2�5� t� 
 ���ERENCE 1��׏7�I�[�m�������2�ԟ���
� �.�@����3ß|� ������į֯�S��4k�$�6�H�Z�l�~������5�̿޿� ��&�8ϣ���4�� zόϞϰ������ϱ�7c��.�@�R�d�v������8�������@����0���9�� l�~��������C��FACTORY DATA\��'��9�K�]�o������ 9������������	 ��GYk
�2_������0���2_� Pbt����' j�?�
//./@/R/ d/'���/�/�/�/ �/�/?'���/H?Z? l?~?�?�?�?'b�7? �?OO&O8OJO\O' 
��?�O�O�O�O�O�O _'�ՇO@_R_d_v_ �_�_�_'Z�/_�_�_ oo0oBoTo���_�o �o�o�o�o�o�o�� /ASew%�����3��%� 7�I�[�m���_�t7 ��Ώ�����(��� ���d�v��������� П;����/��0�B� T�f�x�㟥�/?��Ư د���� ������? \�n���������ȿ3� ��O��(�:�L�^� p�ۿ��'_�Ͼ����� ���߃ϥ��_T�f� xߊߜ߮���_oqo�� ��,�>�P�b�t� ����������� (�:�L����4��� ������������*�p� ��0BTfx�� S����  2D������ ����W��(/ :/L/^/p/�/�/� K��/�/�/??*?<? �/�x?�?�?�?�? �?�?O?�� O2ODO VOhOzO�O�?C��O �O�O�O_"_4_���� j_|_�_�_�_�_�_�_ ��	�o!o3oEoWoio ��o�o�o�d