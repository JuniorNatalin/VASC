��  	��A��*SYST�EM*��V8.2�306 4/2�
 014 A�5  ����A�AVM_WRK_�T  � �$EXPOSUR�E  $CAMCLBDAT@ �$PS_TR�GVT��$X� aHZgDIUSfWgPgRg�LENS_CEN�T_X�YgyO�Rf   $C�MP_GC_�U�TNUMAPRE_MAST_C�� 	�GRV_}M{$NEW���	STAT_R�UNARES_E=R�VTCP6� %aTC32:dXSM�&&�#�END!ORGBK!SM��3!�UPD��ABS�; � P/   $PARA� � �<��ALRM_REC�OV�  � A�LM"ENB���&ON&! MDG�/ 0 $DEBUG1AI"d�R$3AO� TYPsE �9!_IF�� D $ENwABL@$L�T P d�#U�%Kx!;MA�$LI"��
 T�APC�OUPLED�� $!PP_PR�OCES0s!�(1Ns! *�!> Q�� � $SO{FT�T_ID�"�TOTAL_EQfs $0'0NO*2�U SPI_IND�E]?5X�"SCREEN_NAMr {�"SIGNe0��/�+!0PK_F�I� 	$TH{KY�7PANE24� � DUMMYE1d�4d!�54�1�*��ARG�R�� � $T{IT�!$I�� N DdDd D�0DU5�66�67�68�69�70�7G�1EG��1E0G1:G1DG1�NG1XG2cBF�0S�BN_CF>" }8F CNV_J� �; �"L A_CMN�T�$FLAGyS]�CHEC��8 � ELLSETUP 	 P� HOME_IOz0�� %5SMACR=OARREPRJX{0�D+>0�dR{lT(��AUTOBAC�KU�
 ��)DEVIC�3T	Ic0�� 0�#���PBS$INTE�RVALO#ISP�_UNI��P_D�O�V7�YFR_F\0AINz1��1<�S�C_WA�T�Q^-jOFF_� N�wDELZhLOG�R8�1ea�R?�Qf`Ɯ3?�� {1�5�4��MO� ZcE 	D [MZc���awREV�BIL�g?��AXI� �b�R  � O�D7P�a$N�O�@M���cr�"w� Lu<q��`Z0D�C� d E R�D_E�`Ts $�FSSBn&$CH�KBD_SE�UA�G G�0 $SLOT_�V2�q�� Vzd�%��މQ_EDIm  _ � cQG��CPS:`a4%$EyP1T1$OP^0r2dap_OKnr;US�!P_C� �q��T�vU UPLACI�4!TQ?��p( �QC�OMM� e0$D�;�Q�J0f`�y�?�2oh�BL%0OU�r ,K�QQ2QU �B�@y O]Å���CFWt X �$GR� ��M=BZ`NFLI���0UIRE��$g"~� SWITCH���AX_N)PSs"C�F_�G� �� 
$WARNM`"`#!�!�p�@LI��f�NST� CORz-�RFLTR`�/TRAT;PTb�� $ACC�Q��N |��r$ORI��o"�RTlP_SF~g8�CHGz0I��bT�1�uIʐT���K�� x pi#
Qnr�HDR�2QJ; �3I�2D�3D�T F�5D�6D�7D��8D�9�"��CO�D <F ���p��#�܀O_M�~� t 	P�Eq0�1NG�1iBA� Q���q��!�@Qp�0=q�0I�P�P�J�p�G�S���pm �RC �����"J���_R��gC��J�����ļJVep�%C��X���p0푨��AzOF� 0  @F RO��&9�6��IT3c9�NOM_xyV�lS D$��D �0��A�B�'&�EX��B0��P���
$TF��E0��D3N�TO��S3U8P+� N-0P_H�j 1�	E{� %�Y#&�d%�(��1�$�DBG�DE}!_p$Ʀ�PU��1a21)��I"��AX�Ae$�]eTAI�SBUF�iv�Y�/ �� k�f�PI�$U��P��M��M���^���F��SIMQ|� �$KEE:�PAT0�����N#���Y#$�L64FIXb/��⥟TC_��b� ���c��CI�Ύ�PCHOP��ADD��������I"m0p�3�_��!f�� �n!
��a��W���d"�<$�MC�� �0yJBE�ͤz���l�+�i������� ���pCH� EMP��$G�����p_x�lS��1_FPm�8�@��SPE��@lPn�������� V�q0<r�A��JR�<r?SEGFRA��3 ��R�0T_LIN\{sMPVFs!�$�'�_�"�#m�"� �R�$�y� D )���`�����2 �f�)P���Ţq�f�SIZc���T���3�RSINF��G�R �@e3 e��> L�8з�CRC(�AcCCn��3 ���*���1Ma����D��D&�e#
)C+e`TAM ^�&��T(EVT&i�Fj!_
F��N�&�@f�`��((������'��j1���A! 1�>p��-�RGB��"��FB ׂ��De�RN��LEWر�Q�����/�. �R>Wt"� ��Ư��5b�#�R� HA;NC�$LG~��!@�QU�y�gp��6�A:`� a�c�R?2 �3p00��3\��8RAnS�3CAZ��7HP ��O�GFCTC�Y07�F)�p���R�ADI�KO�H@�@�o��D~�.��6�S�p�����qMPW*���M�4AES��l#�B�|���4#  �=I+$�CSX��H�B��$*�?p�s��T�B��C�0N�p�qIMG_HEIGHmq�rSWIDK�qVTt��M��pF_A 8{��B`EXP�A4�N�U�CU7�]�U%�w% $_�TIT���r�s�p��E�:RZ_% {�&*�b{� ��A~�NOwPAD	q?W�i?�,������DBPXW�O�&�'��$SK\���r <�`T�0wTRL%�( �,��A!���@��rDJ���LAY_CAL`�q	��`�@�gPL	�~G�SERVEDW�wb�w��'��	�*��9��0���`AA�%�)�b��PR� 
x�D"���%�g* _���$�{$"��Loy�+|"�,��&�,��"�<�PC%�-��"�8�PENEL���!.�"ќOqsRE}��r/H�0�C�� *$L2�+$os��+@C�T 4�WO�0_D�A��RO�X�X䤍�>|�RIGGE��PAUS��VET�URN���MR_��TU>��a�E�WMF��GNAL����$LA-��n��,$P��-$P\@!�.�b��1C!�!��DO` ���\�H��b�GO_A7WAY8�MOD�0~�B�DCSrp�EVIm� 0 oP $іRB��
�PI���SPO��I_BYT2�����TXw�L$�1 H�� 7��Ф�TOFB��FEl������lw�CU2�DO����0MC��N���7�(`����Hy@W����w �w�ELEGR�3 T����cCINQKh�����U�L��cHA��}$��} pw�����w4 ��`MDL��O 23��(�O��^����C�2����J]�}O�m�}2�U� r�h�������	�����	�w�%U5� $]��0�PcC�PZ� �Pa5бw��ϲ���̵IDJ�˶�b˶W� ���NTV��вVAE��(РW�D�2W���J�&���pSAsFE)���_SV�B�EXCLU�a��N>2ONL���Y6�p�3x@�Qw�I_V�@>�PPLY_���X� Ƕ��_M�"���VRFY_�c��M�S3�PO��x@!֧@1~S4�^�O���İ��@�� 6��`TA�_ ����  �NpW�SG�  7; ��CURπ��}S��tpUQO�REV0�ٯҦ�jPUN�p� �ԥ��Ё�����0����ѧ@��� ����PаI�r8 @b� F���T�OT��At<�At'qAt^� m�`EM��NI�r9 L �`�r�Aʱ��DAY	�LOAD��6tv�Bs=5>q��EF�P$�JX�:�' SO�������`_RTR]QX�; D�!O��RQ{�������:| C7 񙔠�qA;`���< 0��Z��p�Z�>��6DU�5��bCA�� 3=9�[`NSk���ID� PW93U�����V��V_U��< �DIAGr��u>8 *$V��T%ep
Dp}R�r��{V2`7��SWB�� u���B ��;�� �3OH�r�PP2a}IR�Q}B���m�`�����	�BA�����D@������=���CY �RQDMW�MS� AZ`xw0{LIFE�`�/Hq��NB�K@��@��!����C�@+f�NЀY0�AgFLA�4��OV�@�W.`��SUPPIO�`�A���`_���z_X�C�a���Z�W��A��B����CT%U? `>��CACHE�'C"�ۣ�կ���� SUFFI�ϰ�`%a�6t��Bs6>q ���DMSW%U@ �8��KEYIMAG��TMF�C�!с޻&INPU}R ;�G�VIEL �1wA �BGL/�����?� 	tnpfPcBMP�!g1CIN^�Tb��	UBv�JB�a�d��O#QT�3��S��Uu59d�;�|�OF��H���C �Va!gOTF���ץ1�D[�P_GAI�Q���@�@̒��NI_�0C���5��\�6�PTIC��O�P E���"��}1�A{�P�CF�@INy��P[EA�q�@!� ��A|$P�3D  P�*�6D�7I�8T�=ĹRv�=�AVE�FF�BP�c�C���3AW_�@<���E����;DO<4SLO���1TERCE/���D1L/`�J3UFU'RQ��E�e{0�P�E}1�D��B�FE��3N� �3qPQ;`�5�R�6�R^�5��G�FF� 䠣�$�0��G �1�0���1F ����0�3�0 ��AbyB��cCARRg#i0�9T$ <2%cyftqcRD_4�06FSN�p���T� �FSY��D�I"e�C��A�DĔ�dEG�R�F !	Np0u0��Hb�C9 �0ǰY���1�@3��G T2A I� { _��3]6�0��s�1�s�1����D Ц$J�z�STp@!�r)��tk���tv��t���pEMAaI���/1{�SB�@AUL��K�")8}1�COUdP�!|�D9T!���L,�@�2M�SU��ITh�RZ��U'}�N��F SU	BRT��C봅��*r�w�SAV~�@� EAS��m�������P��NM�ORDM�p_RP8d���ډOTT���A���P�60��s��AX��,��XRP�R�'YN_�>�Mb��6$�௕�G3��@;IFO 8���b>=�N� �05м�r�C_RO�IAKO���Ҟ��@R�!8���8��DSP�&��	PA��I(v���ß�R��U���D��M�p�IP0Á��D  >ڔTHRES�`˕2��TZۓHS�bۓR`�E[@��V����@��㑤P��NV��G ����]�ؖRPFB��ad���@(�PSCb�Ru��M-P��FBC3MP�À�ET�a��mO�"FU�DU'���QPPEP���CD�љ[���-3x�� N_OAUTO��P��$z���z���PS*y�CR���C�BE���(v����QH ��в��r�г���@ N����S��k���v���P�����!��7��8���9��B���1�1��1*�17�1D�1�Q�1^�1k�2y�2T��2�2*�27�U2D�2Q�2^�2kʕ3y�3�3��3�*�37�3D�3Q�3�^�3k�4y� ��v�OUT� ��R �� "@	WvPRuPLCWAR+v�`�����R�$FA�Cm�SE��$P/ARM1��2m�"�k��$x³�pA �<�EXT��!S <�)9I�g�0Rv���枵��F�DRdTT @ ����E-�BE8�11(OVM�4T��A\�TROV\�DT��|�MX��vP&8�{���IND��:!
���`E�PG3����� b1�`DR�I�@c�GEAR��1IOQ�KL��N�@:EFF\�k�� |�MZ_MCM1�nEt�F�UR5��U ,��V�? �0@?� Ð0��Ei@� H��p��2� V�RTP~�$VARI�5�̻��UP2_� W *�?�TDI�iA>�TV�� w ��BACG��X T�p@�U�=0�)$PROGC%�?����b�IFI��� wYPa��	�D�FMR2�Y ,�k��B-� Mp�1�8J\s�}0�p�L�_���AC@I�T_[U�C_LM���(DGCLFl����DYt(LD�b��5������4��uZ�!) T�sFS؀�t[ P�P��":2�$EX_�!�(�!1'�נ���!53;56�G����\ ���2��4l�O�N����1�T�1Q�G�R��U��BKUv�O1�� ��PO��9�0$�W5�0�M6`LOO��1S�Mw`E�� �����`_E ] �,0�  �,PM:�5^�9ORIp�1_�9SM_M	�0�`�:A/Ia�5<1U�P:P b� 9-��b]$�5v@�^��G{J� ELT�O�CUS�@ONFIG��A� c1aC�rD_$U+aא�$}��A�@P� OT��G��TAk�-�3SN;STv`PAT`�f`�RPTHJ(�N�Ep� ��W��BARTE` �E�p���r�AR[pRY��SHFTR��AQ>CX_SHOR1�K�J.F 9@$HG�Pa>!�.�OVR����PI�tP;$U�� M�AYLO0�!A��`� ��pQ]���]�ERV� �Q���Z���Gv`QR��0t;e��tRC����ASYMt����AWJ�G����E�?QkibQ�U�d@A�CU�q�P�YUP��Pġ�VO5R@M��?0�1 �c�r�2�6P�@}rs`��q�%d Ƚ��xLTOC�A|�1i$OPo�"����2��pH�O,��Z�REbpRأ��X)�K�ReipRU�u}x[QDe$PW�R$ IM�ubR_Xs8TVIS/@�b*t��B e� $HzC!�ADDR��H�1GR/�$����v�R3�����f H��S��N���\���\���\�*Â�N�����HS[�MN�!g uB�trq�[�OL1��h���^��0ACRO�p�AhqND_C1�|�a�t�šROUP��!r_"ÐI1�Uq"q1��6� 2��<���<�Q�=��`<�*�<�7�6�AC��IO��D7���G�y�� �h $� �Pp_D��0�⣂P�RM_+� ��HTTP_|�H�#�i (��OBJ�E���t$�L�ES��ְjN0\���AB_��T�3�P�S����DBGL�V1�$KRL�yH�ITCOU@�1G�f�LOC�O�TEMPt�����zpv{psSS����HWe�ԫA#�kW��`INgCPU,2�pIO� e���r�����*¿��IBGN�$ql���� WAI�s��aP����R���FW,$ ېLOm��s�|���y�AN�A$Bo��������������RTN/`�CUF_DATA�㖠�����_MG�2/ F�>�S�(SE��r��8REC4���N�bX2�h�}I� m @� �N�_h�Y�3t���E�XEwɒ�Ф d�_�Xu�0�n�$GSCH�`�QP�Rn��FLGvQ 1�	/�oo�����v ���OPÒ�1~�TR1A�B��CS���9�px $C��CTA��'�IGN�MoO҈0�M~�Tֈ��v���vN_PCSO�QUp��ECFBa��Q���u� �Ғ�	\r��L�������@DFRs�������SPT �$���SE3Q_� Z3NS��H� *�ɀ��rC�q�@ Xl�SL�}Pr�Q � -@o�bc��0�se:!���IOLN4q� 8��R�$S�L�$INPU�T_�$�p��P�- ����SL���!r�r��#���ݐF_�AS�"s:$L O$�O��Р�r+�Ռ���PHYP���^� ��8�UOR��#t `J��(�%�s�%�|���pP�s�������|����� T�U�JR�u � rN��UJOG�G�$DI,�$J7��dJ8O	760I��AXj7_LAB�QHpZ �NAPHMI� QY�D� �J7J8�0_K�EY� �K�)�L�%v  �AV8އP�CTReS��FLAG:2*pLG�$w �����Y3?LG_SIZJ��0`>� =A�=FDHI<S�1J;@= :tsC�� �A�pj�@�X_R��x�����5��LNC
H2x����U01#��!BpU�)!(�L�2#("DAUN%EA`�)�Dtd"Z GHEr� ��M�BOO>Q�yt Bd��pIT�Ø${�e�#ү('SCR��`�D��[2�$�MARGI�D��,�X�ct2��M�S�0�L�W�$M�=$X�J{GMC7MNCH�&M�FN�F6Kl7q�j9UFx8�Px8n�x8�HL�9STPx:V`x8àx8� x8RS�9H�`�;U�C�T�3�bX�p7CIU䑌47 �R,6� +�2G\9lPPO�G�:�%�3�d2�OCG�{8���GUIj5I�3�B(3S 43Sh0l1�P�rC9���&�P�!N݁-�ANqAM�Qq�QVAI� ��CLEARfD�n�HId�~Sr�~RO��XO�WSI�W�XS��X8lҸ�i�i1��T�քn�DEV�����!_BUFFqzj� �pT0R$I�EM����'  (
bjqq{� �p���ˁIpOS1je2:je3ja x
b~Q	p| �! ߈�aZSq��{���IDXtAP�ƞ@z�jK�T���Re Y���a {$EvC{T���v)v���ch�} L�s�����������w3��u �Kc�#_ ~ � +�x#��!�s��MC"� �! CLD�P��vUTRQLI � wT2 �y�t�����p�͑�nQD��ڠLp���t�ORG2  B!�'��������r!�|�s͔� �����tE�t�SV_P�T�p��R�ǄφRCLMC݄m�����pMISC�� d%!�aRQ�����DSTB��` 1K��!X�AXvR� |[�t�EXCESm$G`,�M��⡂��?�PvT���㠃�M�_�I�����r����pK�� \�PǻMBۢLICL�B�� QUIRE,CM�O>�ON�DEBU���ML���Ш���e�H�Pށ�p��2�Di �$D�$U�PyACK�ED����DPxv��I-N�b$q�_Q �p \�U�������/��	�=�U�4�T�I���ND:!SSb�#""$f��DC�6$IN]ю3'RSMD ���PNpr�BCs�PST���� 4q�;��fR�Il �e�eANGx�bI���ODAQ��=�;�$ON,"�MFqT��i��00p�uz� 3�SUP�vv/�FX&�IGG�! � �ဃs��#�s6F�tR{�v��b��ɵ��ȵ�����+�D�ATA���ETI�8 ,�+��MH�b�[ t?�MD?�In!A)M���YӇ�U�H#��SX�DIA�Y�ANSWe�Y�Pa�AXՅDl#)8�ŀ���[ ��CUSV��0�I��p��LOf ��������G���5������ ��MRR2>2��� ��J!�Á d$CA�LIQ��GrQD�2�f`RIN�0G�<$RR�SW0������ABCS�D_J2�SEe�I�L�_J3:��
��1SPm I�P����3���ѓ�
I���J����ā�OaIM��CS�KP�z<�- kS<�Jm!�Q<�m�S�m�c���_AZ˂	��E�La���OCMP&����1�� ���`�1���� ��Z��
?��INTEVpSb!���2I�0Vp_N���7�a��3̒�A	DI|�����DH��t6 ���Y`$VQ�l���a$l1$ `�!`��Q�-��2��H �$B�E���	�qACCE�L����� IR�C_R-��ONT<�a�c$PS���rLAp�#�s x-!sPPATH�	�Z�Z3)����_@ga���ʂ�C���� _MG�Q$D�D��"$FW�5�1������D}E�PPABN1ROTSPEE��ka/�pc�kaDEF�ۑ�Ap$USE)_P�>SP�C�@>S�Y
 � ʁ �aYN�1�Ac�x&,�o�x!M�OU�NGtB�O9LJ�$INC�� ����X��'3�Y�ENCSP��I�!�V�IN�bI)52Ќ�c�VE� H�*22�3_U>��<3LOWL�Qz@���p�%\6D]@I�3� �p�%r�C' #6MOS�P��MO���`ʇPE�RCH  y3OV p t"�7�a�3��_2��������b%��P*�A)EL=T*��)�$5p��_:ZFu6TRK�4�bAY��Cܑ�A)��E�C!��`�RTI8���"�`MOM�BX�@ܒc���G��D��C�\jb� DU2��S�_BCKLSH_C)U� �6�0�#���:T�"EZ�!e�CLA�L2`"2���@�`wUC�HK�p�eS� RT	Y���5$�U�0�9_�c�4_UM���Y9C�S�SCL�T# 7LMT��_Lg����T�gE m!`k�P e��0Q�!&@bd&�8PC�1�8H�pl�d��UC뀎rXT� .�CN__�N���f&�SF��9Vb""��7��a)u�hCAT�^SHo�_���& U�Q6��*����3PA�T�"_P�U�C_�p�P�F�0�q�C�t��UJG�����sJ0O�G�g�BTORQU T ��3�I�/��2�A��_W�E�D���7��6��6�I>�I
L�I�F9�)��,#�VC� 0R�J����1����Əc���J�RK�������DBOL_SM�!5BM���_DL�5BGRV�=�6��6���H_p���]d�COSq��@q�LN�������� � �� ��h�Қ����b�Z���6�MY����}�TH��1�TH�ET0e5NK23��[����CB`�C5B�CT�ASƱ��`h������`�SB����k�GTSE�#!C��� ���|s���ϓ$DU�P>G�D��!����3��AQ��&�$NEB��I��#���L$~ O�AS�|���8c�n�n�LPHq�Z�45Z�S��ͳ��ͳϕ@Z�ޖ�����~ V��QV��� ��VźVһUV�V�V��V
�V�H�����µ�:qT��һH�H�H��UH
�H�O��O���OIٴ�OźOһO��O�O��O
�O��FZ��������ԑ��SPBALANC�E�~aLEȠH_S�SP��4���4�>ϖPFULC8�_�G�_�ϕ!
1���U�TO_�P�uT1T2���2N�Quc� ��O�Aa�?�0��A�TK@O���'�IN�SEGu~1REV8B�~01DIFtEF	�1�+�r1�IPO!B!�gQ@��G2�����Q�LCHWAR�
"g"AB�q�E$MECH�� ��!���VAX�APEd��u�� � 
����n5ROB�0CR#B����b ��MS�K_��� P ��_R R���+:!vD1r/0-"+ ,3�ET+ �IN��MTCOM_C��>� �  �3�~ !$NORE3>��OPWO��� ߗ, k SB5U��QOP� ʿT�
U�=PR�UNq�PAR Dp�����0_OU�!��S�AB�"$^ IMAGVQ( �B�P�IM� BI�N'�BRGOVCRD<��	@P!Ap!_��q��R��`RB�`��[aM�C_EDT_� �K`Nl�M�JaPMwY19Ia��n�SL6�" � x �$OVSL��S;DI0DEX�c&H�cKA "V�!$N'! �5 %#:'5(����_� �" � @�@l"���2� �2�
&_���'�!�! ��0�ECT�  ǚ H(��PAT+USP{@CD�Z;DX�&BTM�'�!	I	�4Ia�#�" � D( E"�"�Z�E4��!FILE8J@gP�!EXE� �Q �72K24t#�{ ) �� UPDATZ1$T�HXNDP���x���9��PG7��UB�!����!�!�#JMPWAeI'pP*#�5LO`¤F�p�!�RCVFAIL_C�A��1R�@� �V�a�dx��<E�R_PL�#�DBTB�q�UBW�D.F� U�P/EIGpI��TNL#p�0D�BRT�� ERcVE�c�D�bл1�DEFSP�P � L( ���@``�qp�CUNI"7�@b�1RR0!�.�_L��P�! X�Pr !� 0�q�!N] ATA$�uNP�gKET$R#�BUt�PIPB!� h~�ARSIZEi`�@E0GQ�RS� OR~�#FORMAT���uDCO�Q�EM2���TSUX� :" D�PLIpB~!�  $| �P_SWIp� ����U@p@AL__ � $�AAV�B���CVD	�$EZ1�`C_�zA� � � 1Q�VaJ3��V�80RTIA4hi5�hi6VMOMEN�Ttc�c�c�c�c| B @ADtc�f�c�f�cPU��NR�d�e�c��e�b  �S�P H$PIQ� �6�H�Z�l�~���! ڦ������ ��GQ�&_SPEED�G�R �tE�D�v�DE�,@��v��x��y�ESAM#��F��wL�EMOV_AXI�! �z��%���7�z��@)1d��2dR	 md`��	`a Б�INڌ 	`/����؄B�#�x��#�C�GAMM���A��R��GET�rF�IMS�PDcd
��L'IBR�1�BI�@bS/$HI�0_^� $f��E`ŘA���ӖLW�� ����$� Ӗ?b���@aCfEq��|�  $PGDCK����_.��PdւSiaɅ���c���f��c W�$I� R��DW�0�1"D��LEa�qЫ!�?hᠣVpMS�WFL1DM`SC%R�86�37+�U��qW�4�S]�p7�P��URB����GR��S_SA�VE_D����3NOC`C�!�2Dd���� Sj<v幾Uy�mpʀ���pW�v<Ƚ�.aO�AA��񊅰���e �x��vv��ǜ�Z�\���1�<�QMuߦ � ��YL 5s~�ɇ��~�����N$B�KA���WѰ(��4��`�����M��L�CLK�aDi�^�1j�k��P�M�� � � 9$���$W�Є�NG1]a��d��#d ��*d��1dV@��s��(�S��	`XPO+ca�Z&��P@t� p�| ��Uv������,�;�Ca_�� |�Si���i��c��@�c��mj	���jE@L�� *���y�� �^`��P�Q�PM�4 QUP� � �88PQ�𽡤QT�H� HO��HY�S�PES����UE�r�hP��� � 6B;Q#��#���_� 'Ѵt���EN/	PBG_@B�[ mB?�#*#Jہ���I��pEW �vG�TF-b"�PO>�4�   ���"UN� N� rq�O�rp� PD��E��-3�BROGRA�!�264M �ƗITh@�{ IN;FO�� � ������{ (v�SLEQ�v�6�u6��{ �D$�0p�����Ov���j�#��E��NU�΀AUT���CO�PY���0��qʰM⾑N��^�PRU����� gQRGAD�Jv!�wRX'��B�$P&3�&W(P�(��$�s	 �3EXvF@YC��@!{NS�T� �4A�LGOk�.`NYQ_FREQ��U �w�!�T�LAhC�!��8�b.��5CRE�0��fl�IFQq�NAT��%�$_GhCST#AT�@4��M@R� ��31	���Q31��|$wELE�0 �Nb<�SEASIr1�� �"�a2�1���6Bƀ Ia�"�q��M���2�AB�Q/`E� �pVU1�6BAS9b�5�����U�@� ��$��1F|$��� �X �2 2� 	����QFBPG�Q|р�eE|F �{%PFe1�=GR�ID��SB|P�wT�Ys3p| OTO\ �1Q� �_41!E �BwRO$��$�� ���LI:�P�ORAS�C'v�BSReV0)TVDI�PT_�p6PHT��RW�p�RW4PY5PY6PY7*PY84Q�PFs�e1��� $VALUP�3���4��gF�%�| n5	�b�C
1���0AN����R1Rp�!��TO�TALQ���7cPW�#I�AMdREGENKj`b4�X!G�s�&��fm�TRC�rKaC_S���g``�3V'����c>�1E:3�@��p��cV_H�@�DA}��`pS_YhƱ�&Se�AR}��2�>@CONFIG_SE��`RJ5�_� ��I����D�� 4{�O�v�k�F�sPS��F�f�gC_F��m���!L�����(cMϰ����q�r^⃁z��D�Eհ2�KEEP__HNADD�q!�$�0�CO�0+��A�r%�,�Of�
���q��,�1��,�REMC�+����Bh�����U4e+�HPWDs  q��SBMs!�vB� ,v�cFL�з���YN�p
�M:�C���pQ�Ern�� �l0DB�oMTRI�DA,��B� 0�K�TCLA�����U AYNS9P��֡SEAꠁҖG_P�Tn���Bο�RGIn�QSOCLUK ��P��L)a�$SC`0D�#ےALI�r���S��B#U�A}������� ���w1��_�P�H�TIC�[�`�p[�RE3VIo��OLP����p�FK��_F�SScEGQ���b��;ITc3� �l0C�P��TU� MSEC��MN���̢������`�0�G����20O��1�$N�̡_�e�$�PA� j�P�0vO�iP��MLr Px�� ~�  ������e1��  G$OW-����G�� ��p���Hp2C�Ĺ�Aü�!ߤX�AX0�Q��A7HI��6 ��ٔ�2��Ϛ��2�BV�EP���P�`Q���H�ߢ�r��V�t��`a� B^"$4:�Q������p�M��y�O��l""�SMH��<�M=��2� �L`U_P_DLY��Æ�DELAk�>a2Y�ߔ�� �QS{KI'�� �P��O��NT\P�B��P�����`
��P�� �a��v��l���vP�� �P�ڐP�ڝP�ڪP�ڝ9���J2#����yrEX@T�#z�����z�.@�z������RDCa��� � ��0TO	Rq���	��!�����SDRG��H��k�b��Gg��eER�qUBSPC�G�z�?_2TH2N�!D�~#�1� ���@v��11�� l�p 2�F17��Ta��� Oѯ%��^������SD��VAHOM]E�� `]�2e��k�}��������� +�]�3e������p0B <]�4e��ew����� ]�5e�����*< �]�6e��_q����� B]�7e���� //$/6/
�8e��Y/k/}/�/\�/�/ 8]�Sπ�f��  �AX8^�u`� �]�-ET�yp��m2L.fk3IO�p�:I0  �]�POW>�� � U0K�Θ�]�(d ����2$DSаIOGNAL#gf�CJ���1 �RS23�2q5� ����%8��ICEt�����̳��ITq&aOP�BIT"cFLOWFCpTR003b��UXs�CU+�M�SUXTtđ��I��FAC1D�ų%@ �	@CH�Q� @{p�p��Cf�$�`�`OM,p�_���ETޠ�sUPuD�pA3� �	@�P�@�Q�� !
�(s�A�����)��^.�ERIOc��PT:p3T�2_���Q/P�DAMVWR���/9D���qV��6FRIE3ND(�@�UFi��t8�P���UMYH�p@����GTH_VTE�TIR���R�P~�XUFINV_���ѥ�WAITI����WX���Y7fG27WG1��@1SQbbg2pp_�RE�O_t��s�Q�`��[PC�C�u�Ї_TC3��Ķp�e`��GˀŲtqֱ@ &Q/A�r�jQX�EV��E�a�������D�oX s�ML� ���`��SX��]E#T�C%G3�WCPgws�|t=D�LOCKkuv�`��V��q�ta�$�fB[���pkQe�qY1}X�lP2o[2�{3o[3 }Z�y'�~Y�yC�6.Иs.�r$VV��V8eVl����a�b!�غ��F�sρ��f�qB���`�R�ɠ��E�$߂�S�@a�Tu���PR����uj�qSl�G�� \��B�� ����%s[��w���[���p�@|`��@��
��DS�17� ؚ�R_6�oQ���f0$RUN��A)XSA�`A�PL�QV���THb�J���6��aqTF"�NT���IF_CHeS��~�qU��6��G1��0���ҽ6�_JF�?�PR�`���RT�C� ���GR�Of�A�MBVq̐C�rÃ��`UI#���BU)cRSM}��a`r��_W�P�TBC[_P�PCM��D��ЖLDR��ރ�A衰�@��c�IT�"o ���TA��G� s���|� ��ę��� ���� �ݾ2�  2� ��S��g��	|# �Vд�}�I�t��ˀ~�TOT��~�D|젖�JOGLIzCN
`E_P��qBO���}����`�FK��_M#IR��Ѵ{`M>r�AP]q��E)P�Ҕ�J�SYS�˂J�PG'�BRK�bѕߐ:��I"1  N�pS�Y�x�D�A~��B�SO�}��0N��D�UMMY15U��$SVVpDE_O�PoCSFSPD_�OVRU��� L�D��óOR��� N�P��Fߑ�Ʈ�OV���SFڟ��.�F� �́ճc8ؿQ˂L�CHDLz�REC�OV��[P��W�PM��vձ�ROoC����9_ ��� @�&`�VER��$OFeS&`C;��SWD���r�����Rū�TR��1W1FpE_FD�Oƃ�Ӡ��B��BAL�����1K0%�V�A �B�@��b� �G�,�AM*Ã�D�Z��t�_M0�|B��3��T�$CA���DU����HBK�AЖ��I�OoU��1qPPA�����������2~��DVC_DB)c�0�ё�21���́H�1�P���H�3P���AT�IOˀ�A{���U8tS젆6CAB��nR��c7p���`S��A��_��@ЖSUBCPU�2��Scp�0�B��@�sj�B��2��$HW_C_ dЧs5�sAta���$UN�ITb�\ U AT�TRI�i��CY{CLϳNECA�����FLTR_2_�FI��8���6��Pxǻ��_SCT�cF_UF__�q
�FS�1:�ZCHA��Q�)9�qB(RS�D���2x�ޣ�1�0_TW�PRO����g@KEM*0_��V�T�q� z��D�IPҔRAILAiC>��bMg�LOu��S��9�R܀��䁟�V��PR2�S�a�p�!C$�$@	��FUsNC���RIN�`0Ԥ�'$fARA8 �b� ��P#X0��P#W3AR/���BL�af'$Az+v}(v(DA``�Q!�(�#z%LD�@ ��q�#��Z!ہ�#�TI�5y���$��@RIA�A�2AF
��P;A.3��45�p8�r@�MOI` �ևDF_�P7��Ac�L�M��FA�PHRDYJTORG͢��fS|� �5MULSE�P�����J��J�������FAN_A�LMLVV�AWR=N	EHARDpP�E��Y"2$SHADOWl��/�?Bc�@�w@u�:�_m�ЖAU��`�:�|@O_SBR&�E���JU &�/!��CMPINF��pk�D�!�CREGpUq��л�i�� J�v�Q$;Q$Za��e�O�j��� ��EG�~���*Q#AR�����2�q7Wܧ ,�AXE��ROAB��������R�_�]�w�SY_�dQU��VS��WWRI�P=V5 SCTR����T���EW�8�FT�qkB�`B��P���V,�����OT�O�A8���ARY���3b���B�ƱFI,5�ܳ$��Kq1��JSa]�_�S��EU:3�zbXYZ'B�j�5�fOFF��Rb�zbnh7`B��"`�d��V�  �cFI� ��gq��«�"��_aJ��6���y�$a@ddk6��qTB)qd�2arC� �DU�ҺDV7�TUR@X
3�uAa�BX�P��IwFLg�Tд�7P�p�ex�Z�û� 1�8�K��MДDV����ORQy��V#�W3I��2�+�s0��h�à�Tz�OVE����M� *��C��S ��
R��6@��*A��W  ��<�! �50����� ݀Q�*�������'�S�'���ER��Z!	B�E�PD��e�A����eH%t?g�!���!AX��6��! Ua���˙�1˙�`ʚ �`ʚZpʚ�pʚ��ʚ�ʚ1_�ʖ�0Ǚ�0 י�0癮0���0��0 ��0'��07��0G�d��X�DEBU-$�(!4C����vbAB������~�V��, 
#�Y�?�K�OW� #aW��aW��aW�ZqW� �qW���W��:4fp42\���cLAB�bI�) 6�GRO� Ir-L��B_�L��T�� �`�@ �4�J�0�A<�AND���Z���e]�Ay� ���@~a��0�!�ȡ ~`NT@=!?�SERVE��P�� $�pT Ae�!��PO��K@��-`z��<��_MRAQ_� d � T�Ўe�ERRr2�00T)Y2�I��V�`��N7�TOQ����LhP8���RJ� 0��D@>Q � p 4��Ԯ�_V1f��������2��2���D@��p�H����$WT� ��q�VQ��@C$���d0iӨ���OC�!P�  }�COUNT�Q� h�SHE�LL_CFGQ�� 5!pB_B�ASVCRSR�A)B� ~SSW�!�h�1��%g�2��3���4��5��6��7r��8��[�ROO�0���Y`}`NLQlsAqB�úi�ACK4�IN�T� ���0a@8�0�_PU�0@�OU�3Ps l���I����TPFWD_KAR<ї0�RE�Ę0PO`�! QUEr�t��� �r.@_AI@7�H�{`�8D��EzbSEM?�Ox0)6�TY*�SO��)�DI6�s ��8��b1_TM��''NRQg{`E� (��$KEYSWI�TCH���I��H=EupBEAT�q�E:PLE;��Uҍ�F���SNDO�_HOM20O<#REFe�PR�a���Q�P7�C� O�1�v��O �;rK@0IOC�Mgt��a� �vG�HKQ� Dxa�t�RESUUB��M��"��w�wsFORC�x�#\�G�OM>;P � @�*3*~@U�SP9P1�$�9P3�4� {�S�HDDNP�� �BLO�B  �p�SN�PX_ASP�� �0v�ADD�GA�$SIZVA$VqA:���0TIP��'#�A�� � $c�( �`bR�S��"QC7Л&FRIFHB�S����� NFjODBU��P���%�#�)��  ���Si�P� x6��SIT�TE�sX�.�sSGL#1Tab�p�&��<3íP$0ST�MT�qU3P&P�VByW��%4SHOW]5��ASVDTU�w� ��A00~� �2��7��7��7 ��75�96�97�98
�99�9A�9\P�7� �7ӱ�6�P�7�C�3W�TpH�91�91�91�9U1�91�91I1IU1 I1-I1:I1GIU1TI1aI1nI2�92�9`@X�9�`@X�9@Yp@XI�p@X I2-IU2:I2GI2TI2aI�2nI^�h�93�93��93�93�93�93�I3I3 I3-I3�:I3GI3TI3aI3�nI4�94�94�94��94�94�94�94�I4I4 I4-I4�:I4GI4TI4aI4�nI5�95�95�95��95�95�95�95�I5I5 I5-I5�:I5GI5TI5aI5�nI6�y6�96�96��96�96�96�96�I6I6 I6-I6�:I6GI6TI6aI6�nI7�y7�97�97��97�97�97�97�I7I7 I7-I7�:I7'�7TI7aI7�nD�Г0P� UPDb���"+���
`�0�GUN_C���s `�g�PUT'�cIN\���<AX�|�GO�U
GI~��IO_SCAw�ޒ0YSLOP�� � E%�"#��':' � d�� ʤ	�P��� �R��F��ID_YLj+�HI&�I����LE_g�V����$���SA���� hЂ�E_BL�CK��M1��D_CPU��F ��: &��Y�k�����b�R ;��
PW"���[ 	�LA�2S��h���RJ�FLO 5��5�đ 8�V��|V�� �TBC#��C!�X -$}�LEN��$}��D�RA��d!$��WI_��&�1}�C�2��AM�b��� 3�II�s ]���TOR���}��D����� LACEG��}������ _MA+ �J� �J�GTCVQ�r� �Ts sڒՈ����� �2��JF��$M�ԙ�J���0��� ���2/ ~0���ӱ�JK(�VK:�$�B�3,�J0O�>�J�JF�JJN�AAL�>�t�F�t�n�4o�5��N1�ܥ�d�N�ry�L��{� px��CF/!�T�v�M�?1�"B�NFLI�C�# REQUI;REEBUOy�n��$Tx�2�6��z� �x�. �3� �\rAPPR,�C���{�
��ENs�C�LOS� ��S_Mp� $ ���
�$���A?  �����  ����%���������s�VM_WRK �2 ��� 0  �5��)L �L	#�`������q���_���n�+5UOS<;M_� �����/B/�T/7I�)tG�� k}�5/�/�?� /-?;?1/r?�?g/y/ /�1�?�/�/g?O�/ 8O?Q?_OmOc?�O�O|�I��BSPOSU�� 1��� <�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
���B�~�N�LMT������C  �1�IN�:�L�0�PRE_E�XE]���l�.�A�T}��J����LAR�MRECOV ���l��DLMDG�  "�LM_IF ��d�*�<�N�`�n���������ǯح,� 
�O���FNGT�OL  �K�@A�   4�F���PP<��N ?�������Ha�ndlingTo�ol �� 
V�8.20P/A2�E����
8�8150�������
33713�23��� ��15345����}�����87DE3����	F�.0�14i�FR=L�? 2����:�DX��TIV�}�l�J�i�UTO��� �h�P_C?HGAPON=���h�����L�1	� ��������I���U� 1 ) \����>j� �4����VIQ�c߽߇������ �{��HG�����HTTHKY�� �߬�����6�H�Z�l� ~����������� � �2�D�V�h�z��� ����
������ .@Rdv��� ���*< N`r���/� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ 
??"?4?F?X?j?|? �?�?�?�?�?�?OO O0OBOTOfOxO�O�O �O�O�O�O___,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZlu�*�TO�uχ�DO?_CLEAN��(Ծ�sNM  #���9�K�]�o����_DSPDRYR�&'�HI���@(�� ��%�7�I�[�m���������ǟ$�MAX@Z��t��q���X�t���i�PLUG�G���w�Å�PRC*��B�ϋޏП�?�OD���(�SEGF��K�������'�����%�7�o���LAP̏߮�Ӌ����� ��ӿ���	��-�?��Q�cϨ�TOTAL��0���USENU
̠�� �x���r*��RG_STRIN�G 1��
��M��Se�
~��_ITEM1�  ne��0�B�T� f�xߊߜ߮������� ����,�>�P�b�t��I/O SI�GNAL��T�ryout Mo{de�Inp���Simulate�d�Out���OVERRɀ �= 100�I?n cycl����Prog Ab�or�����St�atus�	Heartbeat��MH Faul<D�M�AlerW��� u��������������� �s���q �hz���� ���
.@R�dv���.WOR�����X�// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>?P?b>PO��8�0 �q?�?�?�?�?�?O O)O;OMO_OqO�O�O��O�O�O�O�O_�2DEV�>,P�?_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o|�o�oPALTD �a��o�o
.@ Rdv����������*�<��oGRI���t��oN��� ����ҏ�����,� >�P�b�t���������Ο��b���RD��� �@�R�d�v������� ��Я�����*�<��N�`�r����PREG�n��0������� �,�>�P�b�tφϘ� �ϼ���������(�~���$ARG_��D ?	����k�� � 	$��	[�]�����^��SBN_CONF�IG kۊ����CII_SAVE  ������^��TCELLSET�UP j�%  ?OME_IO���%MOV_H!�4�:�REP���X�UTOBACK��
��FRA;:\�� �調�'`#������� ���x�1�5/12/03 �07:33:46���ت�B�T���x��숄����������"�����Pbt ���5��� (:�^p�� ��C�� //$/�6/H/'��  ��_���_\ATBCK?CTL.TMw��/��/�/�/�/��INI��`��֞�MESSAG���!��s���|��1ODE_D&���?E_O.P0?��oPAUS�1!�k�� (7�?��տʸ���n==�.ܽ®����)���? 9Ȯ?�?�0I�?O  (On�(O:K$OZO�HO~OlO�O�Ic4m0TSK  s=���M>�/OUPDT'0�'sdP5XIS��?UNT 1k���� � 	 �tE������ q�{ ��C�����GP W�y t`�� ~܆ ~S�3 � � ���8�kU�_�_GPť�t��?D�� �Ӄ^�� �"A�_
��� �ѱ^�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1U@e� v������� ��Q�<�u�`�����ཏ��͏�&TMET�15]Pޏ7�ڏ [�F��j�������ٟ�ğ���!��E���S�CRDCFG 1}k���	�����@�����ȯ گ�����"���E�W� i�{�����
�ÿ.�� ����/�A�SϾ�Y���GR.PPQ?}�j kNAN�j�	��nz�_ED� 1t��� 
 �%-p EDT-k�b��ϼ߻�� @�-(����/����?�\�ϛ� ����2��~a�UP023��&�� 9۹�$�k�d��f��3\� ߩ���
{;R<؅���7�I���m���4(��� ��d���Q�������9���5��d�A����������w��6 �0T���T��C���7���  ��� /gy/�B��8X/��/�?��퀁/�/3/E/�/i/��9$?�/q?�/���M?�?`�/?�?5?��CR�� �<ONO�O�O�?�?�qO�?}���NO_D�EL�ϛ�GE_U�NUSE�ϙ�LA�L_OUT ��  gҜ�WD_ABORT
_{�CP�ITR_RTN � /����CPNO�NSTO��nT ����$CE_O�PTIOkX|�ƣPRIA_I	PRnU�P���PFn��+[ڳ%��Q_P�ARAMGP 1]+[�^g��Qocouo4kCH  ��np�`��`��`��`Ș`ܘ`�  �D�`�`�` *�`*�`4�`>�`�`R�b��`�m��`��`UҘ`�`��`�`e�`�`��D/�`U9�`C�`M�`W�`a/�?��o>ogyT��n|�`��`��`_�� C��p��pU��p��p��`��`U��`��`Ř`ʼpUмpּpܼp�p�`�����| ;Mv��������� �1��ŏ׏���I� [�m����������-� ?�Q�����	��i���PHE�@ONFI�GK_��G_PRIw 1+[ �� ��د���� �2�D��V���KPAUSP�OS 1���S ,]E������ƿ�� �Կ� �
�D�.�Tπz�dϞψϮ���j�O��Q�_�7�QO_�MORGRP 2�l �` 1B��yr�:� 	  :�R�@�v�dߚ߈�k� ������������2�� �h�V��z��:�L� �������
�@�.��Dc�!݋���?o��o��`��0K���1 r����������������PP��+U��` Ua�A-��k}��:
\�	�0P�N@f��5��`�53DB���+YI�2)c?pmidbg[��@m:�� �� ф�UApG�kpE�    -a�E����`��P����-/���0"��0#�g/v/A/ r�0s�fe/�/��|�/?ud1:�/�?�7"DEF Y��7)�!c!buf.txt?�e?4 _L64F�IX , ��?�\�?�?�?�? &OOJO\O;O�O�OqO �O�O�O�O�O�O"_4_�F_~?MC�,P  d�_�_�UfS��t]��T�Ub=����aB�a;�B�� C (B��P�C+�Ch�C��
�;�C���D���9D&�D���D�d�D�F�!mF��fF��0G �F���xG0ٟGt$_�	r�X!���]� �YT_�o�o�o�o�odo vo�o�oO:s^� *���� ��9���s�2g� =S<�	����*����b���ӣ�Sx,�a�p@����p� D*�"�D;πK�3D�m� E�π�@� E��fՎ�`� Eh EE��3F�EZ� F�h��?�  >�33 ;����@s�n,�=�5��=���� A�UL�_�<#�
�2����/����~���Q��̣Q��E��� � #H���-�fJ�L� J�2�Z��J�9�=�e� w���������џ��� B��f�=���a�s��� ������ͯ���� '�t�s�]��ρ��ϥ� ��ɿۿ��5�#�v���2RSMOFST� 6>���9T1>�PDE !=�pcG���;�3��U�O�>TEST�02��R7"�r��|�| C4����
ȹ��!�CzH�Pw��R��s��@i�-J:d�
-�I�_1�#7�-�T_�00PROG %�r�%v?��*�T_I�NUSER  ���(�C��KEY_�TBL  ��(����@0�	
�� �!"#$%&'(�)*+,-./0�12345678�9:;<=>?@�ABC00GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�������������������������������������������������������������������������������͓���������������������������������耇���������������������9�t���LCK���<��STAT`+��_AUTO_DO��%�INDT_7ENB� ���̟�T2�-�STsOP��SXCh�� 2$B� 
 8�
SONY XOC-56L輸��߀@��ʹt( �АOHRC50K��o�7��Aff���// �>/P/+/t/�/ a/�/�/�/�/�/�/?�(??L?^?�TRL���LETE� ~�	T_POPU���-�T_QUIC�KMEN�4SC�RE�0B��kcsc�4��0��9��c_�4U�M�0U 1��_  <K�%k? gOK�EO�O�O/ÁO�O �O�DF<��_�O_P_��LStart �SM Comm �%IBSCMA�NS[_�NEnd�xV�@�U�0�_�]Us�er Cance�l�RUCANCA�C� o�L
�RRe�set�BURES oo3_E_�oYoko��o�o�o�o�o�@Z�ange�GZG_-A�_�ocuL ^��������)� ��_��ZVAG�_KONFIG.�RVW)��=�O�؏�s�-Dateie�L�%DATEI �1�����E��.�@� ��d�v�ß������П�"bMacro S�tep tt�PM�SK_}<��LW�ait Moni�tor3aSHTP �G�L�柫���������ZCYCLE �POW�PPWD������ DOW��%	#�_MAI�Nu�a�%Cb�NUA�L�?�ZCD���&��C�[�	���������?|(��$oDBCO� RI����5#DBLOVR�D�%�NUMLI�M��d���D�BPXWORK 1'���ϩϻ��������DBTB_N1 (7�P�Q����s�DB_AW�AY��GCP� ��=��3�_ALU��?3��Y�5���$�_DBG 1)N�� ,I��
��+(!�Cа�а���>�ӆ�$���5�M�� It�B�@��	�OoNTIM�7����)��
)���M?OTNEND����RECORD 1�/�� �@�� ��]�@��� @,� �x��@�o�G�O逿������?�b���?����RDONE
�TING

 .|�5���#��������� ?����d�������?������@@��@���x�\˴벖���������iEXECU��O"�5)�����/����@� �6���@]Հ@��� �T��@�������^�ٖ���o������]����n�_Qc�����** �c�@����@F� �����@� @?��@��g�g�>r��������� y�BЎ�/�/�q��w��2� ��q�@�-�@�SE ��p@��( @�d�@W����Y��� ���K���������>��� @�O����Ȉ?	0 @����������]~�i����=ċ�f�B�>/ P/�t/_/��/���	 ����/�/b/? ?�/M?�,�"�/�?�? ?�?�?<?�?`?r?'O 9O�?�?oO�?�OOO �O�OrO�O_�O5_�G Q_c_u_�_�O�__�_�>_  CANCELLED
�_o#o �_�_Yo�_}o�_�_�o��o�o:�3�TOLEgREN��B�Bȉ��N�L���CSS�_DEVICE �10�   üƹWi{����������sLS 11,}�K�]��o����������rPARAM 2�����r�r�tRBT� 24,|8��<�I!�D	>� ?��  ���W��K~@�B�۶��D�Ɇĕ�α��{��C�F�B��`OTēA�˖˴�;�C,n�I�C�R�HY���h��U�ő ��p� α\���	����A�Ʌ
��Á�c4�Ɇ���� ������̯ޯ����&�ɍD�DzΒ�j��ѰB�W�A��A���A�A��A���ɊЕ�p��Ĳ�ʳC*�Ɍ��mv�B:�B�33B2p$ffBtff��¿Կ�  uTe Z�� S� D�ɍ)�K�]���E�s� �ϗϩϻ������>� �'�9�K�]�o߼ߓ� �������������#� p�G�Y���»��� �����)��M�8�q� ��^ό�������� ����	 2V h������� 3
i@Rqv ���b�/�/A/ ,/e/P/�/t/�/���� ��/��/�/=??&? s?J?\?n?�?�?�?�? �?�?'O�?O"O4OFO XO�O|O�O�O�O�O�O #_�/G_2_k_V_{_�_ �_�_�_�_�/�O_1o �Oo,o>oPobo�o�o �o�o�o�o�o�o c:L�p��� ���� �M�_��_ ��n�����ˏ��ۏ� �%� o.�@�m�D�V� u�z������ԟ!� ��
�)�.�@�R���v� ��կ����ݯ���� S�*�<���������� �ο��+��;�a� <�j�|��πϒ��϶� ���������]�4�F� ��j�|ߎߠ߲���� ����G��0�B�T�f� x���@��������
� C�.�g�R�����xϦ� ��������Q (:L^p��� ��� $6 �Zl����/ |�%//I/4/F//j/�/�/�/��$DC�S_CFG 5�����!���dMC�:\� L%04d�.CSV�/�#=���A K3CHS0z���/#>^?�?�  ���2�1�?�7�� �`iMU����(RC_OUoT 6�%�!���/�!_FSI� ?I �9#8AOSOeO�O �O�O�O�O�O�O�O_ _+_=_f_a_s_�_�_ �_�_�_�_�_oo>o 9oKo]o�o�o�o�o�o �o�o�o#5^ Yk}����� ���6�1�C�U�~� y�����Ə��ӏ�� 	��-�V�Q�c�u��� ����������.� )�;�M�v�q������� ��˯ݯ���%�N� I�[�m���������޿ ٿ���&�!�3�E�n� i�{ύ϶ϱ������� ����F�A�S�eߎ� �ߛ߭���������� �+�=�f�a�s��� �����������>� 9�K�]����������� ������#5^ Yk}����� ��61CU~ y������/ 	//-/V/Q/c/u/�/ �/�/�/�/�/�/?.? )?;?M?v?q?�?�?�? �?�?�?OOO%ONO IO[OmO�O�O�O�O�O �O�O�O&_!_3_E_n_ i_{_�_�_�_�_�_�_ �_ooFoAoSoeo�o �o�o�o�o�o�o�o +=fas�� �������>� 9�K�]���������Ώ ɏۏ���#�5�^� Y�k�}�������ş� ����6�1�C�U�~� y�����Ư��ӯ�� 	��-�V�Q�c�u��� ����������.� )�;�M�v�qσϕϾ� ���������%�N��I�[�mߖߑߣ��$�DCS_C_FS�O ?������ P �ߣ�����"� 4�]�X�j�|���� ���������5�0�B� T�}�x����������� ��,UPb t������� -(:Lup� �����/ // $/M/H/Z/l/�/�/�/ �/�/�/�/�/%? ?2? D?m?h?z?�?�?�?�? �?�?�?
OOEO@ORO dO�O�O�O�O�O�O�O��O__*_��C_RPI����@_�_�_ �_X_��|_�_o0o+o~��SGN 7���r`�v1���12-JUN-�24 17:14�   ��03�-DEZ-15 O07:3�aC`Ab XJ�a�I,��H���a5n�`wa�������i�ZX�_��o��VERSIO�N jjV�3.3.2�lEF�LOGIC 18~���  	Gh���Ny��]~0rPR�OG_ENB  �5dEs�`~sUL�SE  cu�u�0r_ACCLIM^�v��s��sWRSTJNT�wfra���0qMO�|�a�q/r�INIT� 9=z���� ��vOPT_SL �?	;��
 	�R575@ch�7�4m�6n�7n�50��1��#tNy��*wK�TO  W��o��+vV"�DEX�wd�rbC`)�PATH� AjjA\K�JBVTU211�150R01\ �\  56S\A�RG2\g�m�PA�RADO\�nHC�P_CLNTID� ?vEs �Go ǟ��IAG_�GRP 2>����R�C`
 	� F?h FR݌�Eu  �D�<5l�B�  =�+��B�C�f�T�CVV��C|軑�d � C[m�C@�9kf362 6�78901234�5���  � �;�G�B��Bz�Bߠ�
Q�B��B�A���A��A�
=5j|֠Ba@�  A�`cAp��B�A�C��C��`B45l �5eW�Ba
բ'3�3B#�B���Bߠ��B�ߠo��
=Bz�7�� ��2�7�F�7�U�!��B=qB�R�B�Bp��B���B��
B�RA��Í�����ÿտ[��A�(�A����A��A�Q�A��HA~�wt��6�h��`Q���+�=�O�a�sȓ
=�}���A�\)A���
A�=qA�}�Aup�Am'�eG��Ϸ���P����sɏ��Њ�U����Ѐ��z���s�l��Ae�1�C�U�g�y�[�:���v�'Ў�Ѧ�-�=}�=m�hM��>8Q�U�-�7��8b0u�7�Ŭ}�-�@ʏ�\���p����m@�*�Ah�а��<#{�
��49X=��$��-�;�����5l�Ð�>���C�  <(�U�b� 4����B��S��M�5iA��?5� ���r������:� ������5Yk�M	?+�?G+�����-���GM��G�U�C���P�C`�-��C��X��}�W
���1��n���ɦZH���-��Ҧ�E��  E�p�D	�'��D�ݟ/Ba�8�?W� �?��=�6�����?XF:��CO��p�����V?a��D�*CD�yH/D��tC`���o/��/J�/�"5i�E)�/D��~?��BdG�/? }/&??J?5?G?�?D`����ϧ�?�?�>�? OOD�V��uWO� FO�O�O �rO�O�O�O �O_�O�O_d_v_T_ �_�_6_�_�_�_o�_ *o<o�_Ho"o�o�oto �o�oVoHO: %^I���i�� ��JT%�7:��6� -��og�Iw������� ����	����?�Q� �ox��������ҟ�� �����>�)�b�M� _����������/� �(�ϯL�7�p�[��� ������ȿ�ٿ��� 6�!�Zω?�?�?�ϴ� �?�����+O=O/�A� �oe�w��o��]߿��� ������+���O�a� ?���!�k����� ���'�����]�o�M� ���/���g���G� ��$J5n�W� ���	��"Q� CU7�y���Ϗ� �����-//( f/Q/�/u/�/�/�/�/ �/�/�/,??P?;?t? _?�?�?�?�?���?O �?O:O%O^OIO�O�O �OqO�O�O�O�O_�O _H_wωϛϐ_�_�� �_�_��/o/oo Soeo��9o�o�o�o�o �omoo�o+=a s�o�Y���� ��'��K�]�;��� ���C/�_ޏɏ�� &��J�y3�X���}� ��������-��1� /U�g�y������I� ӯ�ǯ	��ŏB��� f�Q���u�������� Ͽ��,��<�b�M� ��qϪ��?�����ϙ� ��:�%�^�p߂�LU��$DICT_C�ONFIG ?>m��sVzPoegWS�����STBF_TTS�  LT
:����VER��xQ�����MAURS/T  LT�՜ѿMSW_CF��@���ZP��O�CVIEW��A<�����ώ��� ������XR|��#�5� G�Y�k���������� ����x�1CU gy����� ��-?Qcu ������/ �)/;/M/_/q/�//��/�/�/�/�/?��P�M5�B<�xS�� � ���;SCHw 2H<�
�yQ�Schedu�le 1 LW ���R䑏9ZP?)�?M�HA8�1�?zL[A�4>L�Ͳ2 D�?�?�?O"O@OFO XOjO�O�O�O�O�O�O �O�O__0_B_`_f_ x_�_�_�_�_�_�_�_o�TJafeU4ueD5��9*o �9Dz hgno�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x����������ҏ�����5=`6�Jeb�t���@������Ο���	H� V��)�;�M��?�?�� �?u�;oMoo����ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���_o�B�5� G��7�I�[�m�ߑ� �ߵ�����>����!� 3�E�W�i�{���� ����:�����/�A� S�e�w�������S�� #5GYk}��@�I����92�? `�r�c��T����� �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?� ���?����O(O:O LO^OpO�O�O�O�O�O �O�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�&8J \n����� @R#�v��?�?�? H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d��? �o���o�o�o֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tχϘϪ� ����������(�:� L��o���������
� �.�@������ 3. ���6��� ����v�(�:�L�^�p� ��������������  $6HZl~� ������  2D��p�x�ߦ�d� �����/"/4/ F/X/k/|/�/�/�/�/ �/�/�/??0?B?T? g?x?�?�?�?�?�?�? �?OO,O��P�O�O �O�O�O�O_ _f�� b_t_�_�����_��_ z�V�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���PO8�tO�ODO v���������Џ�� ��+�<�N�`�r��� ������̟ޟ��� '�8�J�\�n������� ��ȯگ쯒O0_b�t� ��������ο�F_�_"�4�F���4��_�_ ���_��:�L������ �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ���������^��� 4�F��V�h�z����� ����������. @Rdv���� ���*<N `r�����R� �B/T/f/x/�/�/�/ �/�H�??&?�ϒ� c?��T?�,���?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_>���_ /&/�o(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z���2/ �/��&�8�J�\�n�����/(?ԟ�`�5 n�@?R?C�v?4��_�_ �_h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �_����ԏ揤���� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�򏐟���� *<N`��蟢� � �2�V������ ��(:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? �ϐ�x?�������?�? �?�?�?O"O4OFOXO kO|O�O�O�O�O�O�O �O__0_B_T_g_x_ �_�_�_�_�_�_�_o o,o��p�o�o�o�o �o�o ��bt� �6���� �z?�?V?��,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ��$��?PoX�to�o Do������̯ޯ�� �&�8�K�\�n����� ����ȿڿ����"� 4�G�X�j�|ώϠϲ� ��������ߒo0�� �ߦ߸������� �F �B�T�f������ ��Z�l�6��������� �"�4�F�X�j�|��� ������������ 0BTfx��� ���~�0�T�f� $�Vhz���� ���//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?r��BO TOfOxO�O�O�O�O&� h�__&_�z7��� ��_��t_,��_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|����>�? �O&O�?6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� 2O�O"�4�F�X�j�|� �����O(_����`_ r_Cϖ_4����h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���Я �����į����,� >�P�b�t��������� ������(:L ^p������ � $6HZl �����//*/</ N/`/ƿϢ/�/�/@Z8N_ �2�#?V�?�� ���H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_���_����_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L��p/ԏ� ��
��.�@��/�/�� ���� ??�6?ԟ�_ �_v_��,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $Ͼ_p�Xϔ���d��� �Ϻ���������&� 8�K�\�n߀ߒߤ߶� ���������"�4�G� X�j�|�������� �������P������� �������� f���BTf�*9�/��ҟ� ���Z�l�6��� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/?~�0�8?T� f�$�v?�?�?�?�?�? �?�?OO+O<ONO`O rO�O�O�O�O�O�O�O __'_8_J_\_n_�_ �_�_�_�_�_�_r� boto�o�o�o�o�o�o &h"4F��� �t:?L??��� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ^?o��4o Foo6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬ�Ro�o "�4�F�X�j�|ߎߠ�@H����� �10��k\�� ���ϟ�������� "������j�5�G�Y� ��}������������� B1�Ugy ����������Ͻ� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�߻�O O1OCOUOgOyO�O�� �O�O�OYK�_o�� R_��A_�_e_w_�_ �_�_�_�_*o�_oo ro=oOoao�o�o�o�o �o�o�oJ'9 �]��?�?�?�?�? �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E��?�?�Oͯ ߯���'�9�K��O�{�����a��$DP�M_SIM 2I����ʱt������C&]Y�&U� � �0� DϨ�q���R�C_CFG J�ʵ�!� X�&]���ϸ������� �5�6ᾰSBL_�FAULT K���s�O�GPMSK�  &Tb׾�TD�IAG Lʷ�հSQ��UD�1: 6789012345��xz޻P�����1�C�U� g�y������������	��Y�۽@���RECP�ߪ�
 ��~�ܿ�ߴ������� �� 2DVhz �������9�K��UMP_OPTIcON|�[�TR���}�_�1PMES�;J�UTY_TE�MP  È�g3BȱЅ�A�oUNIT|ׅ���YN_BRK �Mʹg�EDðZE�|�'t�c�x�T�AT��EMGDaI�[��NC#;1Nʻ ��X/K/&^u�&[d���/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>COUOgO yO�I�!�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o�J<OFoXojo|o�O �o�o�o�o�o�o 0BTfx��� ������4o>� P�b�t��o������Ώ �����(�:�L�^� p���������ʟܟ�  ��,��H�Z�l��� |�����Ưد����  �2�D�V�h�z����� ��¿Կ���
�$�6� @�R�d�ϐ��ϬϾ� ��������*�<�N� `�r߄ߖߨߺ����� ����.�8�J�\�n� �ϒ����������� �"�4�F�X�j�|��� ������������&� 0BTf���� ����,> Pbt����� ��/(/:/L/^/ xj/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?/ O2ODOVOp/�/�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_O O*o<oNo `ozO�o�o�o�o�o�o �o&8J\n �������fo o"�4�F�X�ro|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�j�t���������ί ����(�:�L�^� p���������ʿܿ� ���$�6�H�b�X�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� �������� ���.� @���l�v����� ��������*�<�N� `�r������������� ��
�&8Jd�n �������� "4FXj|� �����// 0/B/\f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�? �?�OO(O:OT/FO pO�O�O�O�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�?�_o  o2oLO^Ohozo�o�o �o�o�o�o�o
. @Rdv���� ��_�_��*�<�Vo `�r���������̏ޏ ����&�8�J�\�n� ��������ȟB���� �"�4�N�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�F� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸������  ��$�>�4�Z�l�~� �������������  �2�D�V�h�z����� ����������
�� H�Rdv���� ���*<N `r�������� �//&/@J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?��?�?OO 8/BOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�? �_�_oo0O"oLo^o po�o�o�o�o�o�o�o  $6HZl~ ����_���� (o:oD�V�h�z����� ��ԏ���
��.� @�R�d�v�������� ������2�<�N� `�r���������̯ޯ ���&�8�J�\�n� �������Пڿ��� �*�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ȿ�������"�,�>� P�b�t������� ������(�:�L�^� p��������߮�����  �6HZl~ �������  2DVhz����� �$ENETMODE 1O��  ����������RROR_PR_OG %�%���:/G)%TABLE  �%�/�/��/�'"SEV_N�UM �  ���� !_A�UTO_ENB � %�$_NON�! P���"_  *�20�20%�20�20� +10K?8]?o?4HIS�#����;_ALM 1]Q� ���2<��+p?�?�?O"O�4OFOt?_OUT_�PUT 2R�=�  @ٌ7���$_\�"0  �01���J�TCP_V_ER !�!2/�VO$EXTLOGo_REQ�6�9�SSIZ_TST�K;Y 5�RT�OL  ��Dzޔ2�A T_B�WD�@xP�&�Q-W_�DI�Q S�4�����VST�EP�_�_��POP�_DO]_�FAC�TORY_TUN��7d%iDR_GR�P 1T�  d 	�O|o�m`�YZ:�n��b���m���0�& ����fmc�o�m�dBh��B`�@N��BGpj@<� xP�o�o#I4m��e@d��A�
�=A��G=`��LA"�kt ��g�����
��"g���������<p�P}<��>��<`?�>=(��s��
 G��0  �uAj��U��C�=P��U�@�y��eCߙ  C̖�B�ܞ�x~UUU��UU�\�叀� E��� ��[�P]���P�W�8�M��D@�K�y
ԍ?B�\?Y��`��O\)?E�?�0��ԍ:I���:�o��9q,�(��Ԏ��� ��{��:F��ʙ �Z ~�Ьԏ�o�o00%U6�j	��o0�ۏT�?� x�c�������ү���� ���>��;�t�#� ��9�����ڿſ��� "���X�C�|�gϠ� ���ϯ��������͟ ?������%߇��� ���������,��P� b�M��q��Y���}� �����:�%�^�I� [������������  ��$6!ZE~-� �Q�c�u�s�o  D/hS��� ����
/��./@/ ���v/a/�/�/�/�/ �/�/�/??<?'?`? r?]?�?�?�?�?�?\J�FEATURE �U�U�P	a�Handlin�gTool 'E �pd`�En�glish Di�ctionary�-Av�3CM�ulti Lan�guage (G�RMN) �,�4D St�@ard'F  8�� Analog I/OzG�  ���$�Ag�le Shift�zH��
�@ut�o Softwa�re Updat�e�@}���Cma�tic Back�up+C��4��Aground� Edit @-A��E��@Camer�a�@F�I9@��PnrRndIm��C)E��
Po�mmon cal�ib UI S ��^�MQnQSPM�onitor,B�F�iRtr%@R�eliab�@,B���Dat�a Acquis�oS,B�U��Piagnos�A�A*D�`Zp	�Pocu�ment Vie�we{R.@�@�Pu�al Check Safety[Q� �`!�5Ahanced Us�PsFrP�Q��5@�xt. DIO �kPfi�T `���-bend`Er�rzPL�R  ؂��Ihgs  ,.���Icr�@3` B�WD*D*�� �FCTN Me�nu`v�S^a X}*�`TP In�`�fac�e  ?�9�G Pp �Mask Exc�`_@_`ȁ�@T��`Proxy S�v�T  �t��@igh-Spe�`Ski;T  �;�@�P7`mmuwnic�@ons.@oU��0)qur�`�`�I� LP�A�b�connect �2-A�`capn{cr�`struAB�+C� hK�AREL Cmd}.XG  |���`~�sRun-Ti$`�Env-A4P¤��p�`el +�@s��@S/W-A�i��~Licen�se�S�Vة���pogBook(System)*D���^�PMACR�Os,r/Off{se�@ k4��P�MH7`�@J� �����Q@echSt�op�atpp�R ��Q@iUb�K /���Ay�x`�@��@#X�Q@od��@witchzHG�+(��pR�Q.E�� �@�͆Op{tmڈ,2z͆��`fil�V"��4@τ�@gOw �_��`SB-T�`
S+C�\��PC�M fun�w,B�۱��PPo�TRe�gi�r=p������Pri�PF`� �Щ����@Nu�m Sell�  �0P��"` Agdju-pBU!h��|˕�J �?K���tatu��,B�8�ɗ�Y  �:��RDM �Robot>@sc�oveGA�`�`R�emj�7anqG �T8a9�@�Ser�vo7`��,B��z~�@SNPX b�r�zH�lZ���BL�ibrFC+CU��p�C@ {���  ���`��o�ptޣ`ssagI� ���TCP1 �C8�)E�á���/I�m��d���M�ILIB!�e�U���P Firm�B'G>P	4@�`�b�AccP	UK���EQ�TXJ�-A�;܃��eln8�"�#«���$A4�0�����@Torqu>�@imulayQQ_ ȕz���u���Pa�q'G���I��� P�Qփ&�`ev�. �*�,`USB port SP�iPN`a�P �
��e1�nexce�pt`Y�n�S �&¢1�h'G����VCWQr�8r/rp����d`Vx�P��\� ;�ƾ�� �����S�P CSUI)E�������XC)E���ʄ�Web P9l��e^1�y�O{���/��`d�Qz`�x�p�?�<Z��^Te�Gri�dD�play ��$�e���D.@�W��^e�R��.qJ�$p�`�ԍ�AAV�M-A_�  }qd3epNa�PAxy`,B���\���-A��op�-A��z��Q@-900iA/�350_i�? }�pAscii�a�ΒLoad�P w��a�Uplr�'G� 0P�A���`�opPBA N����A�qW���,B��m^4�CE�`rkJ����¸�CPRU�T���<|PRT/KeybowA�Man^@v���5}!1Qtrl sd��by E-c� b���XMQl:@qQG=uwF G;�`C��P�@_``�%iRs�s@t �t�� ����MQ�prE�s@�f� �@RPyc��@�r��ori` � ~@��DCS� Jo��sc`���^D��a�Blu /� ��PH��<Z� �J�Qmai�n N#ay�.,B���Py����ifi�S ���hDG@�p+Cx��`��Tc�Outp}u�B �h$�-b����imiz�����`YIhAxis|7a�Q �U��h�m��s��  h��� FRL �"`�� ��`�PHMIo Dev�p (���� A@<}qt�eΐV�PM�c�aP̀�b��^�/C֐}o�bL�J���x�o�  FQ<�u��:�P=��d,Ѓ�Q(�8�O���Q9b���lo�Y��o�  (�A�Y�R�OFINET�J ��[��d�D��`�GRAM/J�OG OJ����@��P��@Passwyol�i��K@5!�th��  &��v�SN�`Cli�Q�'G~?,���SP�EED OUTP>�� ���i�`�� ȑ ��b�s�=e����VAG8n�r(Fh���`�!�`vogi 7��B G@�h��#��3zH�@�"��Weav�I�*DCD����V���p<'�6�4MB D <Z�w���i4FROs;w �(pArcҐ�viszS*Di�p�n�Axx�.@Z���{Pell�L^a�;�MVsh�1(F׏���<c݅��p�P�5�@p� �����5ty�@�GP��x����(��#ױ�� � p1`�3ǡ,Bh0��w�./ys��PR ����І�� 2P��Q7� �@@�`MAI9LR��Q�,?`% <�Pu+ ��ל`f�?�x��Pq �n��]hT1G�T��Ф��w40� �� �]!D���s  �i�a`�,�ֳ3o����PT�ᜄp	.�"Dp�S�N`�`cro���M���Re� �p��Syn.(RSS�)  �LU�q�uiry`		 pN���P?����� @��s��s�
�Qest b(0k��m0t-�  )N� �SS��) ՠteHP�3	�FDpS7@��minLj�>0�0Sp�a_�^(ژ.Dp�"r�'�dib� �3k�@���P cR��)�T��Trp�| Xê4�a�a71{apa9��1��Ġ�!{a�Z� t^C$���dspnȴ20�9@`>�!V8.x I�� �&0��#EM�Z$�EQ ñ��3���RFRE+U �e��d%a1�  2��J��s\0� +P��A��}�when arg ��Sp���fi��͡CD�t�i 3U�?*.pc pi�͡�u �� �d R.Skif�W�F,� BCK  a�pAb��v�q�ungP�r����!r��P��!1O` ��I��Q�A F�`b.T�ig/T $J�~Fix up��� l�bof GO� ��QHT'o f��G�p��=mP� ���p�qs�tQ�P���9��-PS-s�rPI��X��Diff.�a.d S.PN:�FW-CHK ���P���J��}CD:��S�STEP̢BWD�P(R�P��.Er�.af� 8xV�ag_C. 3�,1��sseJ�� �Iss8` �����+P.Alloc.Mem.�~�  �� ���~�� I ���|Q쐀w .K[�l V�ar.Scr �� J����F�B_CMB�lar�����h� ��I�w�r.�!FUNC-?M �Ї�U�-��\��	s �K��Q�˓�"n.sMP D Z�cmd.er.-P�dl.�Pr h�s����c����#rignǱ�& ���j��ATSHE�LL Hepbe�at� ډ~3�No�.On�/��w.SRVO �V��p���,�9�m�� aw����=X GunM.�DO.@!.Gen=.�A ذ�\����?�.scrn f�reeze 7��W�P381�+Inv9`ig.���chP;�d�>Łx ABC&"g�P���,�'!.d���.uP�p.��a�r �_n��4�.��.abd PGPX  :�:i�.��spddѐ�4� ��J �<ځ��4�r7��۳�/H�տ��@8��Û<�<�/����)�K��:�c�E�gè��daσ÷y��<}ϟ�`���ϻ���+е������x�����a�<����H>�	߫��+r`%�G�H�Cy0A�cӿ�r!]ߞә��yߛ������߸�<N<����|OH�������^A2�߫Ąy�'�+a!�C�8�8=�_��6_Y�{���9�u��O��|ϳ�����������������<���L�2B�#����p�@��<�[��B��U�L���(q���*� y����d|)�����Iq�X�����`p���.@���^};��~�.5W�}Gy�Qs|k9mΏ,�}����s���\"��K�3��2�sv�ԗp����1G��<Mo��'�i���~ ���s�ءc^������_�o����#���</3#�U-/O#Ol�&�I/m%���$F��]�/�#38��լrh�$��d/�$ढy�/3�
>�?�o�ҩ�Ϛ����E?g3��טσ4�}�/�4�S��?�3�ϕ`��4q��E�?�W�<�?CJ��	O+C��,��%OGC��y�/cD? �]O�CB)��?�D�0�}G�O�C��1��O�C�F�?�Dzg����O��\OZ%|
!_���p=_�_Sew_lY_{S5g$s�u_�4�K���Ő�t_�T�X]�P��8~��5.4���#d^2��?dgz�z9o�D��?�wd��̔O�d0�s��o�c�0�t���d�żD��dcP��os1�P<�os^QkT��j5Ws�A���Q#$�p�_,3"e�SDWh��~�(��o�tDp���sk��X�զ9p���,^1�S���~qM��d�:��������V�����U:�o߄�� �ُ������؏�eW���3���uH/O�u�PǜI�S�>�+e�����{8�����wdA�pof�� $�V�� y՟��P.U���~*��3� ���)�K�h:� �g�3~_L����������w����s�۵�Kd9c?ѯrb oFt|	��+��R��%^��lc���\����p_�O���` �����h�~���� sTͿ4;����3��'�](3P�!ϧ��r4_��X.�{���o�f*A�ϗf1�$��Ĺ���Ď�4D:����G@9K�#���O?���
9$O"%D�[<U�w�/cpiqߓ��_p->�߯�CP��H�ߺ�9 ���63�J8o��� <_������;�$U3w�5��$���s��L �Ϗ�p�WyY���VT�����^QS�����;9?xO��
�0v�g���+t��4�S�t�<M�o�9s(?�eU�߅����T������$�9�,���4V�ߪ6sk���?$|�KdG�-O�3�_I����̿E��������9֝������ts����|�2tϞ# ����9��>���EKds �T߃;$P�o�u�"5�C��=<����@�p���4AH�_$��T9�	/�1%/Kds�N��c$RtWp��z�I�\/�$w�|���aX��$n�s(r�/�#� �fN���/RE�?�C4�߄�/_4y�0�{4����u?�$�H�n%���̭?�ݰ�nE� ���?s�<�x�#D��\�O?C>��X?�u��/uB�=qO�d?��}v:�(��D�Fp���Dy�y2�O�d9,h��O �"B_;S�s��D�k�Q_�sS�@;�m_�S@� ��_�SQf�<��T�����_fes�V�_�SvS��d���P�7d`�y �Sd�$��MoN?�Zio��e\�J��o��s*�o�c�z��&eo�R�osb sѻ4t	��-�Os�K��Iks�s_�Lo�t�p�_�.E}JJ��s��9�0o�t�
�?Z��;�o�!Uk���T�bpO�����E�Cd TO"u�y�lA��M���C�T�]�����<?󄸰(����.�	�+���,�%�G�{�"�U9!�F�f�;y����<��D�����Ay���ӓ�$z�͟��䰔���1y��'����!��g�'@���x�<Y�{��W �u���ό�����$��Ϥ��8O�ussW����}����#�w���f�O�̔�Be��(w�z�9������ �Zugdh$��+T�c��:�p���Í<����H5�52?�8 �2]1ߠf�x�3"��&PL�R7�8"��C8�0�  S�>�J614  �a�X9ATUP�? �Y�545�  ^��;Y�6�  �P��VCAM�`;)��CRI�����~��UIF�����p�628  �w׌��NRES0�p��A�63.�Vwp��A�SCH�@���JDOCV  �(�����CSU  B��u�Y�0^�ta@��EIOC; ���A�54"�� ��z��9�� ����SET  ��^v��J5�����(��J7�������MASK  �t��PRX�Y@����7 � �2��OCO  ��0�1�3  H��q"��1�R���@���Q����vq�39s�@h�����H�L�CHN��A=�OPLG  ��#���J50~�Jw��CI�HCR��ށI�CSj�����<�50�����`�J55^�����I�DSW  ���[�q����B���q�_��D�I�PRr� d�{<��fд�~��R�o��A U�CM��Ϙ�@P1�^���s�6��fА��xӞv����1�f�l��F��v�� ����PRS*и���QY�9z��$�FRD��C H�bA�MCNS� ��f�93R�J��p�SNBA���\����HLB  �� ۉ��M���� �����(�zq�2R���B��TCj������TMIL?���v��78��,����TPA� 0�vA�TXG`P��)�{EL��ҡ���^��}蠝Y�8E������A�.��a��aY�95����TЋ�fгK�UECN� 0�f���FR��R��`��C������VCO������L�VIP.�辱݃��SUI�@̸uY��X�9W���WEBj����ú�Tj���P�R{62���Q����G�4B��IG���¬^�% PG�S�`����IRC�.��~|�s��·p��89v�8w���U��,L�nX�ð��H6���T��A��ҴsV�y�ֱTL�ܳ���(�R6���L�[���0��Uq��-����v�!��1q�7�R��߸�R53�^�����J68^^�u�����6~�w�<�R74���7�`��~Ъ�s�\	�v���@�wJ56��U)D�]5���7%� 0@�A���@[�`��J98v���q���f���` �J82�������1Ҳ���A�56���P2HЫ .���:Ϭ�5~�_��_=�6R���x������Aމ�6�����\���v�ϛ ���.��Js༱����p�]4.��~���J������9��l�s�p���^h(�s�.�r� ���~��������Ѧ�sxH��^���\_��`(��6ǯ�  �в�������~А���<�҂�}����^��F"�����R��06^��0{y���"0����v� ` SVMr��š��LIrЁ?������dP���C{MS��|k�"�j��q���TY�.���ܩ^�p���t��TOj���$\����T�by]9��@�`Y�NN���o1K0f�o8c�L��RS�ЯB�@���8R�p� Erq�.�cp��i�XT6  ���� F��f���O�PI6 }�2 S�ENDڱ��!!{B�T CPRQ_���L����z��Sd2���0�2�fБ���TSn6 ��@��LM*��  �`�i�J0*6��52^�*�� ���(�<�TOAv�q=��TRAN�o����VA��w}kR��IPN.������H@.����`��EZE�0r���UPD~��:�� 0PMC~БH��P1I� ΀��E0����|�Bv�?���Л@����0}�B^��0�8���@��k�(�B����8@�A�:��,S�B.��� ܙBf��X�RT2v�2���@������@��lm�`0P2QA�e<�A�ѥ�5R�A�z1��P~С���X�P2}���)Q2n�����L�P2���!}��sP.���s �5R~Т�,L �sP��ࠐ$�P24^���p�7P^�ׁ� pR4�����!��3U�w��@P27�����8���P��r���7P�����,pQ3���� A�U�4�1���p�U�5�}���aiQ�Q���P�5Iᐭ�AP33�~�����������=e`T���=e�}\P=e� {��=e2f�`=e�F���=eƿ�xf��(=e�ﻰ�=ehv1`f���������P��� J=e] ��=e(8� =e {_�=e���2=e��P�f0%t�f"��=e����v0*r=e���=e�a��������f8V�f0����=eX,��=e�$�=e���Jv<�� ���{1�=e�+t�=e��=e�dZ�ߝfF��=e��?�v8���f�-��1-v$F0=e��$��=e͏�$n]v�@��K�v� �6�f�`��=e�����f��&=e�\2�=eH����v�T�v��mPv����f�{��v��|Ӆf��F��v���f�{o��f˙a�=e��V�=eX*������f��p�ҠW=e>B{ �=e��,=e����3=e ���f��,vp�vްv;� ]=ey�{@7=e@�A��fwz ���Y\=e��M�Z̗n�fC0�1�A�d��+ `f�`�}�=e�0��=e� ����7Pv���̖��==e������f�F�vw1\=eP�̖wd[v���v�K ��������=ea <��=e��ቆ���=e���v{w�f�|�w��f���醷 >��r�l�א��	v��w����v�<����^Pvo�o=e����Y=e.X���=e"x\�fUgޘvt0�q��4���7���(�޴��(ѾA��=e=�	V=e[w�>�=e���l�/�࠽����e�D�Pv���v�w|@=ew�;�g�,	`f�� 趜�"�=e:�|�=eۃ��f&S�<=eCTlh������t�=e�w@��=e�.�f�؁�v����=e_TDv����4��� T���m�=e,
k��K�o�UHU������� �U�G��w~��=e�\H�����ƚ�����f@|�P�u����vɲ�
nM�kWiu� ��o@X�z)�؟�v�B�؍���Q�=e��x�)� t�f�R�f�?�af�~~�=e�=���=e�:})��;��v�p�w�� �E���t�y���Uf��M�n�=e4�$\v�����	v�`f4P�f=e���Dv��ݍt����xƕs���	v�����Z{6=e^@9=e����I�Lt"�=eJ\!Ϲ橷�^�����=ev"{�9=eZ� #�{�߰�� ��=e��=e+ �ޠ�o��1�T@����^�̖[���;=eպP�=e}{kĶ�/�v�Ȧ���*�<=e����=eŷս����I� ���.~�%=eL��x�^���|����یZ���0��f���=eڷ;UvZ�̖�&QH�J D�f^��=e{ ]�v�9�x<�|��8�����9*�v��=e	}�����0���8��f�@��%]���fG��v6$>v��h�y����(�Em�{��=e@�8��7�s=e�B�`f��U���:�݃����`fʡ�p�fH�?=e$����=e��;'�@�(��|��}lc��P��|�7`�E�:�|����� �<:��� 8�v��&1��X�f^{Q|8 ��)��v��(�vQ���Hfbfa=eл �v �<&Q���<�$�H�{���f�h�醷0p�e����f�w`�-����f���P�pΐ����@v1��0�(�8�4�f*aĶ���D�^�� � �b��P,�>��H55�@Ya�4vA!IP��:!Ip#d.!IXw��@!I�na0J�RBy!I��^�!I �`�!I��� �!IQ��!I��!I��{�!I��b!Iʠ!I�JD��J��!I��{�!I:� �J�	3!I&��!I�!I{�{"!I��!I﫨��JI4F�!Iъ 8!I�J� `JX�u
!I�{���JyBp!I�L��s!I���P!Ilp�!I��!؊!I �W�!IH��!I唽0�Z�`9L!I0��? !I^���!I��@Zt��0!I��Vk�Js{��!I3
��!I���j@ �N�!I� �j� kސj�!R!I��� J��]0J���TAj,8�!I$�RKaJ��KV���qJFA�!I�{�@`Z�x,QZ{  �Z	�f�!I�?2�z1���!I���!I= ��!I�׾�J�w �1J�	!I��,*!I
����A�pH!I/:{A>!I��?!I�T`30J�U��!I�@ h�J��ހz����!I��{9�!I4#�o!j���!I�)DB!I,�(�a!I�A���!Ie��`Z�z@�!Ix`�)!IO��O!Ii���!I�@$�!I�ý��J�2��1j%��J$��!Iaw
P_!I�QR@�s`�$���Xj�RP��J 9@z�jX���3pz{��Z(�J�X�|!IoX({v���DЪ"��zwh��z �0Z�<��z���!IqΤ�Z�^��!I8�#!I �"�@��E- ��{o�ZqV�!Iw|�w��eZ`���Z�!I>�V�`��q��Azz��`�������9:��j�\@j���`��r�!I��۷�aJH�pz�W�{,@� {���nqjh(�J
1���=@��JE>p���@J!I��`ޠ���rp!I� �(��J :Y!IU�;/�!I��³�Jh�zkt�!I�B�!I� ��k�|���V���~� ��c{ �Z��Z�Tcޠ��ߜ١z�L횱j ��j4f�I!Iu0�Z�������Z�J���Z8��j�ݠ�ʡ��j����j��!I�w@��J ���wѬz� �!I�(��z��y'�:�W�!��4^!����!��!�k�� �!� A���!�p4{@!�	
�H�q��!�!�O��^�!��v�!���;&������!��:cP!���:)�!���p�!���� 
�9���!�@U<!���@F!�>���!�����!�� {~�!�)� �!�y�� !�`�!�P}q����!�����"��⑽�!�8����z{ �!��Cţ!��|`�
����!�P8�!�3{~�!���2!��b7�
@�>��&���X��@X����(ޡ���}��{� T�_��Q���aHޡ8:��Г�� *�@$��*�`� ��&�ޡ�jgk��c���j��@���z����`ޡ�})�PJ{���$�k��Q~ˡ��P�W� �; ޡ�k�-�l�{�r��l�d��e��ڡ��<�0:���*����{��t�R�� J�r8��ޡ�<���A{ ������⾡�@H���2p���Ġ��ʸ�
^����?[`�A*d@J���;ޡ:����:�S�!��?L��{0J�������+̠J��ޡ�r:�����ߡ^�� *0w8��� �0J�� ��:ዱOޡ�:ม��쿰2Y}k�*q4���>�,��w�VAJ� ��J��<�����J��`:��.���)0:��8��J0:�.� J8[�>AZc������#J���QZ��0:;�� 0:O@ZJ�y�Z������s��"�q�ģ��*�@-]��*r��eK��������@zo�N�����0�QZp*����%!*�=��w����J2,�*�T��zQ~����x�j:F��Q*Ő���A������*k���~Z���{��:� �!jwT��*��U!Z� F�A.�z�{�|@z�LHQ:{�?�:���	�� �5Z( �ޡ"D���,&ݑ�:�� :�>{4D��,�q*�!��j��j,wz�wAZW��J���P�D��onA��J�1*H�z�TZ��*�;���p!� :�lݲ��r21�@�ޡ���A�?�J���p���Pݿ���`z �_��� �J��9�JrPz���,�z B0:ޅ�� jrm(��J���h�j�\�:�Sݫ�J1I���{�á[��w(~�Кʀ ������A j8�����Z� ��wT8���`�!����&QJ| �J�p�V�>�.�v�j� z����>`D�zY���Q�ܒ$�*ѯ^�ӧ��JN��ݪ�$;�����>�J�*��88�l0:  �?A�� j4��Pz�ݭ�*1*�����Z�@?0:����j�RQj�{�������<<\� ��& 4`J" ��<a� p�Z& �L��*��0�Zq������Z��� z ���ZR���К�cx�{{X$��,�B���d >�������*���ev�J@@J,�P�w���0:x�`0zw(�`�*@ؐP*�������2���2M��z5�6�1ZaP� *�x���=�������E���ߐ������Zh*� �� ��a�p`�V��dК,�1����=@ʱ�@�����u�{��	����zl�7 D�pj��(��:^�B�~����{K @�o(fqz�Zf��*w`�zc�J�*4������0��*� 0�0{<��J�iNA��T�Pzb�T�Z���K�S0z�${ނ�~�o��r��J`��o����1����Jo�fA���0j���.�P����X� �J�A� A����@���0Z�E���������6@��{B�`�@��!J�A�+c`�C�G���S�Jw�ʱ�sѹ1Z9��Jy��P��� � ���0jH���]w ,��|)J�|�P}'��} X j(ف�����g �`�STDz�]��LANGk��{�Y1E )� %E�`P�%E k�%E@�l%E����%E���%E=`(%EAf{��%E�;�%E�,��%E�,�p%E� r}%E8�� %E�!��%E΢�%E�λ �%E��F��P0/%E	�in�F� aF�Fo �VUFJ�HF� ��%E$}�<%E�^K&%Ep���%E~)}_�%E���%E� {
v%E 8��%E�� r"�V�`�%E�^�!%E$���IG}k%E»%�%E���,Vw�"�FhP�F{*?HF�H�%Eo�;��V �HF�(��HFAh�:�%E�=��Vt;��W`�HFH@�0�%E�jHFBX���V�BUFT�A%E,�i�%E'�\|	%EȀ��%E� ��F3Q;��%E�GPJ%E�{^g v��8�%Ew�`Fq��HFo���UF:�HF�ٞ�%E��ސF��%E���SlF����%Ew	�VfMf{8�F��$%E�_`
�V۰��%E�(@ft��%E�H �F:{��%E��;vw̝.�F��a%E��Z��w ��F �H8�V����RBT��p��]�{��@_��d�x�`_�� ��OPTN+����H���{ ������W��t��ލ��0@����:Ȇ��~ō�d�,����:�[ ލ�x�uD��b��|��l{4���w���������o�|���Ѝ���3Q�"��5�W�����������ڢ;ލ�}p?}{�[��ʀ��o Po���P�Pގ��­_���\�������@����0���$�9΍���0@�����Ŗ�5f���{�|Ж��8����#��"����������3{�H�)?;1���^?p0��̔3^T��2K�a�`���}J�D{PN)@>@�����%&B����
�:����8��A��}w��p��k̞Ȁη�B� <���� �<2��	� d{j̵�|����L]�x����ס��!� ����{�h���8y���������/0�޵��� ص��S{0R���Db4���z�Hn��r������4#���`�������*X�ᶀ����2����HK���07)~޵�"�����？h$�����*��aY@���K��(��@��C;USy������g���ߴ�g�ۜ��e�, �g�;k���g��@��g�l��Be�kg�e�x =�e�yRP�g�@�*Ve�灙t�g���e�K �ešs�VX�gì��@��g��z�4�g�%$;�e�ņ�g��؁y�e�0w���g���"e�`s$���g����v��8x�}":���g�9�e�HP{K}e�Xab�e����ke����ͺ�ְJ�o� ��Pe��p|�P{}�e�;�,e���9��g�����e�bÜ�������9X �E�����E�H{E�HViE��X]�GQ� ���E�P��E��A{��E�q�LE��H
$E傠@��E���qE�Tw�(E�a~������kE��@��E��ű E����;E�A���E���"�����E�@��(� {cZE���E��V�E�,����E�����E�BwZ]}�$��E��U4���+��E��������ý�E咷��E�����E�����E���'E���VE悆�E�hw�Q���R�E����"p�`]��v�����������*6�B $��}���E�xB�xE�ZaF�����&�`$]h�$�E�D�����~�Q�D�P� {��P构rd��w�a�E��r:p��(�a�E�Cq~�CE���
-E屷ޒ7�*Pt�Bwxhz��"�E��w�@Q����E�p��E������F�FE�~��Z��a���w���E��"1��E�0��9_h����b��a)��.��E�|��E�w�N!E�ā�P�wu"��&�@��"��E��� ���h�gjE����|=QK'M�
�Tq�Z-�]栦�' |�.�\��u���_E�X�$�E�9 P��8;h
���Ԙ���x?�PRE�o��h��s�~]���E�Q��`D�w?B��]E��w<��(��E�(f=$��$Qf��)&|�������0-|M��`��7����] �� �'$H�'�@��T��E�[�� X�Ehp�&�{R���U�PE��c�a���UvQ�Wv&f��,d)E�G`W��:�E� �0��6�spE��{A}�^���&{a�P�o�Kq��o ��=<�{B�P��}6�?�E�u������f����q������E�n�$�@V �|��ߠ�t�� ������q1
� ��@V}cY��U!��F�����]*�6���}&)3�v�pD�Z�z(Vw�R|�� `��oP=E�;��Ww���V�A��w}k�F�>�twdz�0�@�<wWj�潣+V�A������An�P����~���o,�/�A&��Fw��j�V�U��w��4�&*�$��w�?�,�<&�<�B<��7.{�&�PrE���`G��.ѡvE�L��(��x7w���E�z�0�w���f4>���o�a���&�dF�\��`E��Pޠ�H5�����b�&��^�l6HR��r�Ľ�E� $:�6���&�^)�ϻ�E��������062�D�����V��ߤV���@V��ԈE�$����V�P�6$��&VP$nE�w*�,9��?�����V��&��q��q��QL�Z���(V@8��v���v޾����LPd&��Tt���t���v�;8������o���E�t0�w�f���t;#LV�H�O6�ߌv���4��@�6���4PFU��v8 �d&�@��q���������E樻C9E����2�<6��W�b�k��&��(�E�»+��&�� LV\���L�¿�L�0��'�f�����4��v�Q����x�b��v��,�9F��<�������{�(V�V��F�r��v!�  �
V���� !�G�N����F����F��� �,g9�F(Rs�	�F����� �&�_�}JJv|��h�`99���	,�$FEAT�_DEMO U����3�;� cp��N�D�Vσ� zόϹϰ��������� ��I�@�R��v߈� �߬߾��������� E�<�N�{�r���� ��������
��A�8� J�w�n����������� ����=4Fs j|������ 90Bofx �������/ 5/,/>/k/b/t/�/�/ �/�/�/�/�/?1?(? :?g?^?p?�?�?�?�? �?�?�? O-O$O6OcO ZOlO�O�O�O�O�O�O �O�O)_ _2___V_h_ �_�_�_�_�_�_�_�_ %oo.o[oRodo�o�o �o�o�o�o�o�o! *WN`���� ������&�S� J�\�����������ȏ ����"�O�F�X� ��|�������ğޟ� ���K�B�T���x� ��������گ��� �G�>�P�}�t����� ����ֿ����C� :�L�y�pςϯϦϸ� ����	� ��?�6�H� u�l�~߫ߢߴ����� ����;�2�D�q�h� z����������� 
�7�.�@�m�d�v��� ������������3 *<i`r��� ����/&8 e\n����� ���+/"/4/a/X/ j/�/�/�/�/�/�/�/ �/'??0?]?T?f?�? �?�?�?�?�?�?�?#O O,OYOPObO�O�O�O �O�O�O�O�O__(_ U_L_^_�_�_�_�_�_ �_�_�_oo$oQoHo Zo�o~o�o�o�o�o�o �o MDV� z������� 
��I�@�R��v��� ����ُЏ���� E�<�N�{�r������� ՟̟ޟ���A�8� J�w�n�������ѯȯ گ����=�4�F�s� j�|�����ͿĿֿ� ���9�0�B�o�f�x� �Ϝ������������ 5�,�>�k�b�tߎߘ� �߼��������1�(� :�g�^�p������ ������ �-�$�6�c� Z�l������������� ����) 2_Vh �������� %.[Rd~� ������!// */W/N/`/z/�/�/�/ �/�/�/�/??&?S? J?\?v?�?�?�?�?�? �?�?OO"OOOFOXO rO|O�O�O�O�O�O�O ___K_B_T_n_x_ �_�_�_�_�_�_oo oGo>oPojoto�o�o �o�o�o�oC :Lfp���� ��	� ��?�6�H� b�l�������ϏƏ؏ ����;�2�D�^�h� ������˟ԟ��� 
�7�.�@�Z�d����� ��ǯ��Я�����3� *�<�V�`�������ÿ ��̿����/�&�8� R�\ωπϒϿ϶��� ������+�"�4�N�X� ��|ߎ߻߲������� ��'��0�J�T��x� ������������#� �,�F�P�}�t����� ����������( BLyp���� ���$>H ul~����� �// /:/D/q/h/ z/�/�/�/�/�/�/? 
??6?@?m?d?v?�? �?�?�?�?�?OO2M  )HHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t������� ��ο����(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ������0�   1�,�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&�
8�:�-�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO�&O8I�$FEAT�_DEMOIN [ ;D�h@�4@}PDINDEX]K�lA�P@ILEC�OMP V�;���AkBKE��@SETUP2 �W�E�B��  N �A�C_A�P2BCK 1X��I  �)�MAKRO900�.TP:G_4@%�E_?Z&_c_:G�E1__UT1]_C_�_D�_y\2�_�_UT2�_�_1onoy\3ooUT3eoKo�o�oyU9H�lJ4@�@8u �(��^�� �)��M��q���� ��6�ˏZ�ď���%� ��6�[�������� D�ٟh������3� W��P������@�¯ �v����/�A�Яe� ������*���N��r� ܿϨ�=�̿N�s�� ��&ϻ���\��π�� '߶�K���o���hߥ� 4���X����ߎ�#�� G�Y���}����B� ��f������1��K�@�P�O 2�@*�.VR:���RP*�����#S����yUn�P�C��RQFR6:D��4��X��T|@ |�y�_@I�xV*.Fq�%Q	�<�`�STM ���" ��RPiPe�ndant Pa'nel��H�/��/�Pi/�
GIFs/�/��/F/X/�/�
JPG�/!?�?0�/�/q?��JS{?�?�RP73�?O?%
J�avaScript�?�/CS�?(O��O�? %Cas�cading S�tyle She�etsTO~P
AR�GNAME.DT�O�l�\�OUO�1��D�O�O	PANE3L1�O2_%�_[_��_2P_�_EW �_a_s_oZ3�_:o@EW(o�_�_�oZ4Xo��oEW�oio{o�D�SHELLp�A %+rCm���G�ZG_MENUE0-O�u�q��~�EEINGAB�J�%3�K�L������vSUMM_VA'G.D>?�O:���������yTPE_STAT:��;�S��y����UIO_S3ET�o֟%�A����o��$��yVWEMZROUC�U�C�[��������;�AGV�UPK�]�ǥ߯���0���E;�INS.XM�[ҏ�@K���aCu�stom Too�lbar���yPA?SSWORD���?FRS:\Ͽ��� %Passw�ord Conf�igόG�CONF1����AS�����ϣyEXTSERVOϯ������ �@���d�߈ߚ�� ��M����߃���<� N���r���%���� [�����&���J��� n������3�����i� ����"��/X��| ��A�e� �0�Tf�� �=��s/�,/ >/�b/��/�/'/�/ K/�/�/�/?�/:?�/ G?p?�/�?#?�?�?Y? �?}?O$O�?HO�?lO ~OO�O1O�OUO�O�O �O _�OD_V_�Oz_	_ �_�_?_�_c_�_
o�_ .o�_Ro�__o�oo�o ;o�o�oqo�o*< �o`�o��%�I �m���8��\� n����!���ȏW���{��"��$FIL�E_Dɡ 1X������� ( �)
�SUMMARY.sDG#�۝MD:W������Diag� Summaryx��=���SLOG���p���۟���0�s?ole lo5ϣ�	TPACCN��v�%^�����TP� Account�in=���v�6:I�PKDMP.ZI	Pϯ��
� ������Exceptio�n$�ի��MEMCHECK���������/�Memory� Data����� �)��HADOW������)ϸ��Shadow Changes,��ߴ�K�)	FTAP���χϲ�1��mment TB�D��ܷ\+�)�ETHERNET���͎f���3ߪ�E�thernet ~3�figuraC������DCSVRF�ϊϜϵ߸�%�z� verify� all��cĐc=xu�DIFF�ߓ߸��:ﹰ%��d�iff<���f�z�CHGD11��*��� Q�����7��}�2����C� q��j���GD39�8 �2��� Y����}�UPDATE�S. ��ЋFR�S:\L��U�pdates L�istL͛PSRBWLD.CM{�ό7�N0�PS�_ROBOWEL��g�:SMp�)���M��/Ema�il��aïcį����Տ���� / ��$/�H/Z/�~// �/�/C/�/g/�/?�/ 2?�/V?�/c?�??�? ??�?�?u?
O�?.O@O �?dO�?�O�O)O�OMO �OqO�O_�O<_�O`_ r__�_%_�_�_[_�_ _o&o�_Jo�_no�_ {o�o3o�oWo�o�o�o "�oFX�o|� �A�e���0� �T��x������=� ҏ�s����,�>�͏ b�񏆟�����K��� o�����:�ɟ^�p� ����#���ʯY��}� ����H�ׯl����� ��1�ƿU������ � ��D�V��z�	Ϟ�-� ����c��χ��.߽� R���v߈�߬�;�������$FILE_�7 PRF �����������MDONLY �1X��� 
 �q�H��l��y� ��k���U������ � ��D�V���z�	����� ?���c�����.�� R��v��;� �q�*<�` ����I�m //�8/�\/n/� �/!/�/�/W/�/{/?�/?F?��VISB�CK#��2�*.�VDM?�?0FR�:\f0ION\DOATA\�?*20�Vision VD file�? �/OO3?AO+?eO�? vO�O*O�ONO�O�O�O _�O=_�O�Os__�_ �_d_�_\_�_�_o'o �_Ko�_oo�oo�o4o �oXojo�o�o#5�o Y�o}��B� f���1��U��������MR2_G�RP 1Y��C4  B�s��	 .�ҏ�πE��� �����πP]��P�W�&��M�D.�K�y�
�?B�\?Y���N�O\)?E��?0���:I��:�ov��9q,(~��A��  ����BH̃Cߙ  C�ȓB��З��zr�D	��C���@UUU�UU���S�>�w��j����:
����9�~�:I�;EdlZ���~� ���ܯ� �9�n�Ə d��D���������� οϊ���:���_�� ��nπϹϤ������ ��%��5�[�F��j� �ߎ���J�\��߀�!� ��E�0�U�{�f��"� ��F���������A� ,�e�P�u��������� ������+(a �߂�d���� �'������� ������� #//G/2/k/V/h/�/��/�/�/�/��_CF�G Z��T ��/5?G?Y?��NO� ����F174606 �  m�,��RM_�CHKTYP  �0�s���00���1OM�0_MIN\�0r����0��]X��SSB3[�� �
ADe; C)O8K���TP_DEF_O/W  n���PGIRCOM�0aO���UNC_SETU/P  ��%O�O��O�O��GENOV_RD_DO�6}��mEUTHR�6 dzUdT_ENB�O{ PRAVC��u\�7�0 �� �_�/�_�_|O�_� �_(o�_Lo^o �_mooo�oyo�o�o �o�o$�oHZ�o~���3ydQO�@1-b��s��eB>�8�?��<�
��;�.���3��.��'�˭�N�3G�Q�`���)ٚ��Ȑ*�0��x��g7���B���r�	�y���!�&���"�D�F�x��������l�ɏ������1\�>��:� \�^�����˯Ɵ����ܯ ��At�V�'� R�t�v���ѿ�ޯ�����OGRSMTkScrY�p�0��m����$HOSTC2�1d�y�0� � ESTb|U@ hare  Q�S�q�����172.26.1_8.230����obback\�� 3�E�W�i�Qߑߣ���������~�	cfg_fanuc����.�@�R�b��SH�AREgwPC �S�Ε���� ��r��/������1� |���Z�l�~�������� eVWUSER us������e�� 	=��eB ���mۉ��� �s۩"4FX{�|��anonymo������+y Oa:/u�Q/�/�/ �/�/�/�/ ??$? G/��l?~?�?�?�? �/#/�?7? Ok/DO VOhOzO�O�/�O�O�O �O	O
_U?._@_R_d_ v_�?�?�?�?�O�_-O oo*o<oNo�Oro�o �o�o�o�__)_ &8�_�o�_�_��o �_�����[o4� F�X�j�|���o�oď ֏����Wi{%� ��x��������ҟ� /���,�>�a�b������������ίCʏ�E�NT 1e���  P!a�����	�F�5�j�-���Q� ��u�������Ͽ0� �T��x�;Ϝ�_�q� �ϕ��Ϲ����>�� �t�7ߘ�[߼���� ������:���^�!� ��E��i����� � ��$���H��l�/�A����e���������Q�UICC0����!�172.26.�18.841 G#���	2�s���!ROUT3ER��!7`~��PCJOG7�!192.�168.0.10�CAMPRT�c5 x1����RT ��%/�N�AME !��!�KJBVTU2�11150R01?RS--KU1��S_CFG 1d��� ��Auto-sta�rted2�FTP=��!T�V��/�� ??1?C?U?��y?�? �?�?�/�?f?�?	OO -O?O��/�/�/�O�? �/�O�O�O __�?6_ H_Z_l_~_�O#_�_�_��_�_�_o�o 	SM<����O�_to �O�o�o�o�o�o�_ (:Loo�o��0������ �2� D��ZC��og�y��� ����Z�ӏ���	�,� -���Q�c�u�����TH C����'�I��4� F�X�j�5�������į ֯��{���0�B�T� f���ß՟��ҿ� ����,�>�	�b�t� �Ϙϻ���O������ �(�s��������ϔ� ߿�������� ���$� 6�H�Z�l����� ������5ߛ�Y�k�D� ��[����������� ����
.Q���d�v����4(_ERR fF*���PDUSIZ  �] ^w���>~WRD ?�%�:��  �backup��  uest�gWi{��6#�SCDMNGRPw 2g�%� ��:�] kD@K�� 	P01.�03 8�   �  S ��[  ( � 9� ����&��������������?������+-,�UQ,� 	 � �k@
b+/��� P�; �? .; ���[��S/� � _  N�p��I{/� ? d; ��������O���/�!5U�0�,��d/�!/3/E/2���1?234567&�? ��?�?�?O�?*OO NO9O^O�OoO�O#;�O �O�O�Oy?�?�?F_�O V_|_g_�_�_�_�_�_ �_o�_	oBo�Ofo%o �o__)_;_�o{o �o,)bM�q ���Io���(���_GROU�h*�	-0P	�!�1�cz���B�QU#PD� 6��C����TYP�� T�TP_AUTH �1i� <!iPendan�������!KAREL:*$�-�?��KCT�d�v�L��VISION SCETM�ԟ��]J� �ٟ�I�'��?�9����]�o��������C?TRL j����
 5�?FFF9E3ȯ8��FRS:DEF�AULT2�F�ANUC Web Server2�
�,>۬����Ŀ�ֿ����WR_C�ONFIG k�� f2��IB�GN_CFG il��2] @] o<#�
~�BH|�C��@4:�~�L�DEV�`��V�>� IO ma�I��EXDAT n|����EXFLG����T�FIL o�����O�TP p�Yݮa?���������	MERCA�TOR!RECO|�� "R_ACH60^��ISTW*�V��,�V� "SENS�P��TXQ��99F1	Ke�ine 0�k �h�]%IBSC�����M�4�8�@�E�W�𛩀�T�LM�TN  ���� ��������x�l�X�SBAD��z 7�^�xT��DL_CPU_P5CQ�]B�B���� @�S�^�MI�Nd� =��RT�GN��O�H����рINPT_SI/M_DO������TPMODNTO�L�� ��_PRT�Y����Q�OLNK 1q�@9K�]o���MA�STE����SL?AVE r�b��OZ���UOހ<�CYCLu�$��K�_ASG 1sY� ����aП՗�~���`�%0c�������a�� ����%/0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b?pt?�?�XNUM��z��IPCH?���O_RTRY_CCNQ�I�D�N؁��8�� �Zt��FO�T�S;DT��OLC������$J23_DSP_ENB�0��ь@OBPROqC�C���	JOGI��1ukL�ad8��?����O�??"�ۯ4_�pQJ_o_ �_�_R_�_�_�_�_�zO�y8!�O-oo )_;_�_�o�o�o�o�o��o&oJ�B1 +oeNaoso�o�� ���(�:�L�^�9���BAc������ ���*�<���`�r� ����q����C����?��BPOSF�OF�K_ANJI_� K��&�RE_�.Av/���/�����KCL_�L��2�?�EYL_OGGIN7��������$LA�NGUAGE �����ENGL�ISH ١�LG�-Bw �T���T�xJ ����B����T��'� ���Z��MC:\RSCH\00\Xﶠ��?ISP x���0��⍊�ߡOC����Dz���AݣOGBOOK yY�$�챟X x�	��!�]�x���``͛ўśه	ε���>��ϼ̲_B�UFF 1z(A�ϟ��ߞ /� �K�]ߊ߁ߓ��߷� ��������,�#�5�G��Y��}�����DC�S |ؽ =��͑�L���$�6��H�Z���IO 1}"cJO��(����� ����������#3 EWk{���� ���/Cn��ER_ITMhNd ��������/ /,/>/P/b/t/�/�/ �/�/�/�/�/?��q�SEVڐ�mTYPhN�l?~?�?=��RS�0����B�FL 1~|�@��OO(O:OLO^OLpO�?TP��y[2}��NGNAM]���6ˢ��UPSc�G�I�0c����A_�LOADPROG� %�%UP�054}O��MAXUALRM�ܑ���筥
DR�A_P�R�Dܐ³ڑDPCf�ع�ͪ_$�;Y��P_GRP 2���[ �T�2T�	Z[1\0�P;�_ ���R#oo oYoK�Go �oso�o�o�o�o�o �o*<`K�g y������� 8�#�\�?�Q���}��� ��ڏ�Ϗ���4�� )�j�U���y���ğ�� �ӟ���B�-�f� Q�����������ǯ ٯ��>�)�b�t�W� �����������ݿ� �:�L�/�p�[ϔ�=W�D_LDXDIS�A�@+;l�MEMO�_AP�@E ?�K
 T���� ��&�8�J�\�n�DP�ISC 1��M� �ϻ��T�Q���߅�� ��2��V�h���w�K� ���������
���� ��R�d�O���o���-����������*��C�_MSTR ��,=ISCD 1��͠���� ��:%^I �m����� / �$//H/3/l/W/i/ �/�/�/�/�/�/?�/ ?D?/?h?S?�?w?�? �?�?�?�?
O�?.OO RO=OvOaO�O�O�O�O �O�O�O__<_'_9_ r_]_�_�_�_�_�_�_ �_o�_8o#o\oGo�o�ko�o:MKCFG� �X�ogL_TARM_�b�Xw�b �c��� (t�b_GRP?_DO �X�a�����L��uq?k������o$MMET�PU��Xs��`	N�DSP_CMNTp��`�Q  �I���q�al�v��PO�SCF"��f��R�PM!���STOL� 1�X 4@�`<#�
���a��  �����"�d�F� X���|���П��ğ� ���<��0�r�\���SING_CHK�  %�$MOD�AQ�c��o?�i~��DEV 	X
�	MC:C��HOSIZE�͛`Ȭ�TASK %X
�%$123456�789 M�_���T�RIG 1���lX%�ܪ��c��Կ�� ��˿Ͽ�<����7� ��+Ϩϋ�aϣ��ϗ�0�����/�YP����`��EM_IN�F 1�w� `)AT?&FV0E0%ߜ��)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ������H�����D���AL�t�/������ ����߸����� M� �q������Z��� ������%����[ � �2����h�� ����3�W>{ �@�dv��/ �//f@/e/�/D/ �/�/�/�/��?� ��a?s?&/�?�/�? v?�/�?�?O�?9OKO �/oO"?4?F?X?�O|? �O�O6O#_�?G__X_�}_d_�_�nONIT�OR=�G ?�� �  	EXESC1�c�R2�X3�XE4�X5�Xp��V7�X8�X9�c�RkBOd �ROd�ROdbOdbOd bOd%bOd1bOd=bOdTIbOc2Vh2bh2nhU2zh2�h2�h2�hU2�h2�h2�h3Vh�3bh3�R��R_G�RP_SV 1��q� (d�?��Կʸ���n==�.ܽ®��Ze��_�������Y7�_�D@R���PL_N�AME !>��Y��!Defa�ult Pers�onality �(from FD�) �TRR2hq �1�����Y�  	 d���ŏ׏��� ��1�C�U�g�y��� ������ӟ���	��,�2��K�]�o�����@����ɯۯ��<:� �)�;�M�_�q�����@����˿ݿ���"�
�;��P*�g� yϋϝϯ��������� 	��-�?�Q�c�u�D� Vϫ߽��������� )�;�M�_�q���� ��ߚ�����%�7� I�[�m����������������� E��� E� FZ��|�<N�d�tl~c���! ��   ~q��'EK i�������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? -�F?X?j?|?�?�?�? �?�?�?�?�O0OBO TOfOxO�O�O�O�O�O�O�M �_$�=_�� a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �oP_�o�o�o�o�o�o #5GYk}� ����o���� 1�C�U�g�y������� ��ӏ���	��-�8 N�\���j���� � ����r �B�8� f�\�n����˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�>?W�i�{ύϟ� ����������O�/� A�S�e�w߉ߛ߭߿� ������ _�$_=�O� �s��������� ����'�9�K�]�o� ����b���������� #5GYk}� ������� 1CUgy��� ����	//֟8� N/\����/���/�/ȟ ڟ7/?��??&?8? V?\?z?���/�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_>�W_i_{_�_�_ �_�_�_�_�_�R_/o AoSoeowo�o�o�o�o �o�o�o ��+6�O �s������ ���'�9�K�]�o� ����b��ɏۏ��� �#�5�G�Y�k�}��� ����şן������ 1�C�U�g�y������� ��ӯ���	���/8/ J/`�n/���/|����/ 2��/ψ?�?�?2�8��J�x�nϜϩ��$M�RR_GRP 1_���������  `��X�, ���~�� @D�  ��?�����?������@=�N�Ũ���*��;�	l�	 � ����X��'���F���^������ ��k���K�s�K���yґ&9K�?�MK2�d�s�A�S��߈��?�f��?�;g������Ѡ߯��I�ۿ��6���������X���4  ���  �o����7���A����_�ߏ��s����B�������������(�(Ѽ����  �����>��  ���������	'� �� )�I� ��  ����:��ÈM�È=��9�e���@u�{� v������������Fv����@�?�?�@&�)���C6�B:�BB�C�B�B��Q���^��C��[�2 �		`	`��*��ȕ [; O �	B�� ����Dz��O��$J!�B@e2�j Xy��:y��? ?�ffؿ�<�O ���,68��/(*	ѝ�=$0(��V%P_(z��xU�UԿ�>�33��5;��;���y�"��$;�UU;�ҍ��/�A0�+����� �?fff?��?&�0��@�|g@�;��2�,%5� q1�-��]?��|? �'A���?�?�?�?�? �?OOAOSO>OwO�F5F� fO�ObO�O N?�Or9�O+_�OO_:_ s_^_�_�_�_�_�_�_ �_o o9o$o��lo2o�o�O�oXH(��G�-�G�4��������?EJ,�C'o $6�*p7���~`r����BH�o���o�����qA� A��t<�	��� �w���;��s�(�R��� �d����l���Ĝ��Ç��{C����@ CZu ��c~��&~��~�0��DBTZC5��BjZBa:^�B8�@����%���33��C�C׼���
<#�
?��%�H޸���
��z�BO�_��V{}��%��@�ffB233���B_����L��d��%�L��J�;��I"�PI?���IU߅F�k��ў��5K���I��PH�H��I"��F�B����TK�,k�J��I:��Ie-Gv�l ��Z��W�����w���<����BZ2-��ǯ�����BV�-;����yR<4�?�H��\�g��J��r����J�A�i��������� �=�(�a�s�^ϗς� �Ϧ�������� �9� $�]�H�)�d�oߨߓ��92zu��t�����h�8��&���ƸT�6�G @�o�u��&�"<���LK0�����LM�Z�J\�����8�#�\�G�l� ��}������������� "XC|g����(�3p$�S��!���3GK���s��<-273a��M_����3j��B�}����$3�����@�	/�-/,V�P�"	P_.Z�{o�/��/ �/�/�/�/?�/*??P8:\�F?s�s�wa? #?�?�?�?�?�?�/mo 'OOKO9OoO]O�O�O�J��O�O    XX5�O
_�O_�@_._d_Z52 E��� Ezs�En�WFZ�fB��p,�q�C���pn� ��_�_�_	on�1oP?�Sf�Qf�Y|o��o�o�o!��P�af�4̱s��14�0�\;
 �o,>P bt����������:T�JfXsMtX4��T"A�O @D��V�?�>]� � `?"�-d�A�XU�U?f;��	la�\!}�ો��e��0F��a�������� '��0}�G���?}�h� ����ş��V������0V_�z&'��9�G�8��k��+UUp�s�=��ͭ���Y�s�0�ۯ�Z�&f����G�TY3��u0  '�@[�e�Z�������  ���ҿ��B�P�� @n�.čRCp!��Tϛ�x�cϜ�ćυ�k`����  �kb:v�a�`x#a����
�߮� R�dۖ�8k`z߈�>Ρ+`i��������F�>Ls� ���Aso ���4��e�G�a��*�?fff?-�?&g��σ�&ib�-mv� ]���[���L桄x�� ��5� �Y�D�}�h���p������"o F�P ����7��X��* �&������ �-Q<u`� �����N/r ;/�_/q/�/�/4�/ �/V/�/�/?�/7?"?�R�_4�P�Qp?/? �?:(�0�~?�?�?O �? O9O$O]OHO�OlO �O�O�O�O�O�O�O#_ _G_2_k_V_h_�_�_ �_�_�_�_o�_1oCo .ogoRo�ovo�o�o�o �o�o	�o-Q< u`������ ���;�&�8�q�\� ��������ݏȏ�� ��7�"�[�F��j��� ����ٟğ���!�� E�0�i�{�f�����ï ���ү����A�,� e�P���t�����ѿ㿠ο��+��(�����M�_�I��m� �ϑ��ϵ�������!� �E�3�i�Wߍ�{ܶ5%P%�P����4� ��B����	�B�-�f� Q��u�������� ���,��P��߹�� ��������������� B0Rxf�8���  2K�� *<N`r���������/"/A�F/T*
  T/O7�ߓ/�/�/�/�/ �/�/?#?5?G?Y?k?|��t/��{J��4Ӏ� ���1 @oD�  �1?��3 � `?@��2@��A�X�5���? �;�	l�2��}��KC�0"K> F�ê��?/.�?:&� uO�L> �8�ObO@/�O �O_�O%_]�0@J_`XW�x_��AЙ_p�X_�_U+UU�_�_=���okiS`/`�09oGh�R&f]o�om�2�	�o6^u0  '�o�h�_�o_�x,�2ZO2�hB <Px~ @@��u@�EC���o��o�����R@�&�4��  �@�:h&Nq�~U�2�|j�|��C �в�ċ�q8@�ڏ�>.a�0�1�z2�$�L�">L7a��pA�=���;���@��2��3�2�p?fff?�p?&ǐ��?� �2�4�y�5��8=� ��D؟q�\������� ��ݯȯ����7��@�Ffp&�s�"��� ���2���뿆���� 3��W�B�Tύ�xϱ� ����������~_,��� S߮�t�ҿ��߿��� ���ߔ�
���O�:�s�^���AfpA����������� ���o��?�*�c�N�`� �������������� );&_J�n� �����% I4mX���� ���/�3//0/ i/T/�/x/�/�/�/�/ �/?�//??S?>?w? b?�?�?�?�?�?�?�? OO=O(OaOsO^O�O �O�O�O�O�O_�O _ 9_$_]_H_�_l_�_�_ �_�_�_�_�_#ooGo 2okoVoho�o�o�o�o �o�o�o1C.g�R���(������{����� '��7�9�K���o���@��ɏ���ی�P��	P�Y��~O��x T�~�i�����Ɵ��� ՟����D�/�h�S� ��w���W���=�� � �6�$�Z�H�~�l� ������ؿƿ��� �.�  2��T�f�x� �ϜϮ����������C�(�:�L�^�p߂�8���ߴ�
 �ߓ� ������)�;�M�_� q�������������{J������� @D��  �?�� �� `?��!��A�X��I� ;�s	l!��}�k��e�%�����F���0K����������� ��=�����=(a L�p�y���������z�+v+UU03=���m�����&f�������u0  '/'(K/vo/��0.���/Z(B �/�.� @\ �%\!EC0�_/?[/8?#?\?�G?EP0�?�7  %�P2:�֮!
�!��W<�?�?n? �O$KV18P0:OHJ>��)�M:�?�O�/���>L��V0A�@�O�?�O�?P3!��|!�� ?fff?� ?&'PR?C_O4.�"Q .�M9�}_��_Va� 8_�_�_�_�_oo=o�(oaoso^o�oR]�`F� �o�o�o�on_ �Y�oK�ooZ�~ �������5�  �Y�D����R��� ԏ2��n��1�C�U� �Oj�|������ӟ��l���A� A���'�0��T�?��E� >�����ï������� ��A�,�e�P����� �������ο��+� �(�a�Lυ�pϩϔ� �ϸ������'��K� 6�o�Zߓ�~ߐ��ߴ� �������5� �Y�k� V��z��������� ����1��U�@�y�d� �������������� ?*cN`�� �����); &_J�n��� ��/�%//I/4/ m/X/�/�/�/�/�/�/z�'(y����? ;	???-?c?Q?�?u? �?�?�?�?�?O�?)OPOMO;Lv�P�BPN��{��/�O8�O�O �O_�O&__J_5_n_ Y_k_�_�_�_�_�_�_ o�Oy�Co��LoNo`o �o�o�o�o�o�o�o�8&\J�jw  2o�����@� �2�D�V�d�� ��������Џ�o��
 ��]OS� e�w���������џ������+�{B4����{J��$MSK�CFMAP  �-�� �wvD�E�  ]�ONREL  qE�t�jp]�EXC/FENB��
r���ο�FNCƯ��JO�GOVLIM��dt����d]�KEY�����_PANp��-�)�]�RUN���]�SFSP�DTY�@Ȧ����S�IGN����T1M�OT���]�_C�E_GRP 1�-�t�\��	�� -�?ϗOc��sϙ�P� ��t϶��Ϫ��)�� M��q߃�jߧ�^߱� ��������7���[��P��H��l�]�Q?Z_EDIT��n����TCOM_CF/G 1�j����)�;�
��_ARC�_âqE�UAP�_CPL_�դNO�CHECK ?j� pE��� �������� 2D Vhz�������NO_WAIT_�L����װNUM_?RSPACEg�wr�=�7A�$ODR�DSP^�ѨOF�FSET_CAR8����tDIS�r�PEN_FILE���=���SPTION_IO#�5���M_PRG %�#%$*/".�W�ORK ��$��hpG@S% �mD�C���m ��m!	 ���m!<�����TRG_D?SBL  -����z��/��ORIE�NTTO����Cٴ��s�A rUT�_SIM_D��q�D�TVXLCT� �#B�@-5_�PEXE�g6RA�Ts0	�ѥi4yUOP �<>%�.����?�?�?OI�$�PARAM2೏����>&3	 d��VO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_���_�_ o#o5oGoYoko}o�o��<�_�o�o�o�o &8J\n��@^"�o�����P� 
��.�@�R�d�v��� ������Џ���� ��N�`�r������� ��̟ޟ���&�8� J�\�+�=�������ȯ گ����"�4�F�X� j�|�����������C�߿�3��� !��D�R�ĽĽ���p�� �ǰϦϸ��� �����.�DO]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� �����_������1� C�U�g�y������o�� ������	-?Q cu���#��� �x�	-?Qc u������� //)/�M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m?</�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�Ol� ο��O4�_(�_P_ ^��O�ϛ_�0���_ �_�_oo2oH�aoso �o�o�o�o�o�o�o '9K]o�� �����Vo��#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y��������� �x?ޟ�-�?�Q�c� u���������ϯ�� ��)���
�_�q��� ������˿ݿ��� %�7�I�[�m�<�N��� �����������!�3� E�W�i�{ߍߟ߱ߤ_ ���O��_F_,�:_P� ^_�߂_��_<o��� �������"�Hoa�s� �������������� '9K]o�� ������# 5GYk}���� ����//1/C/ U/g/y/�/�/���̟ �/�/��?-???Q?c? u?�?�?�?�?�?�?�? OO)O;O
?_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__NO�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o ~�����F�,:�$ bp��o��0�B��������D� ��$PARAM_G�ROUP 1��gX���L�`L�X�, ��q��� @D�  &��?�����?�p��F�qC*�����t��  ;�	l��	�  ����X�΀π퀯�^������� ���pH�kI�H�ز ��""�H�	�HGww��|�#�o�oi���qB_�  B���Ҏ�������s�4  ���  �o�������������ȟ�s�BH'���.���q�h���r ,�2���G��sωρc�~�|�  ����������  �Д�����u	'�� � ТI�� �  ��l�=��������@�"����F�ķ���P�w�����������CݐB�B
�C�B��б��Ŀ�ֿ�  ^�C|��@�	`	`3�*A��<�[� ��M�9BUȷ� 3�t��qDz������Ϧ�8����ȦB@�٩0� �;�;�:˅�!�D� ?�ff�{R�d��� ���ߪ���8�����ڰ�HD�����(����P��!�A�����f�>�3�3D���;��;���yL⏸$;?�UU;飑�6��� A0s봂�����q�?fff?�3�?&����@�|�g@������,����©ᵄ�ɤ� ���#���脃�X�C� |�g������������� ��0T?x�� ��q�m�� >);t_�� ����}�/�:/ �[/��/��/�/�/��/{�pސ/�}�2����BH�/3?�/�W?B?g?�?x1AM�A�4㠰1�?;�y7��Ju�?y3o�Ϗq<?�?�@I�Or?�OO:ObEĜ3�Ç�^OC����@ C@5�OO#%@��%@�%O�CBDBTZC5��BjZBa:�^B8�@����`M��33��C�C׼���
<#�
?��̞H޸���
��z�BO��V{$P��`M@�ffB23�3��B_�����L��d��`ML��J��;�I"�PI?�ؒIU߅F��k�x^��5K���I��PH��H�I"��F��B�_�TK�,�kJ��I:���Ie-Gv�l`Oo�O�W�A3oo8WoBo�Z2-cono����o�oBV�-;�o�o��yR<�o�oH���J��r+6J�S^���B�O ������>�)� b�M���q��������� ˏ���A��O�:����!5�����g�h�8��͟@��Ƹ�oݟG @����&:�<F�A�LK0�K�V��LM�ٽ{�EqJ\�����߯ʯ��� 9�$�]�H���l����� ɿ��ƿ���#��G��2�k�V�(d�3p$�S{�4�����d�3GK��Ϯ�_����<��Z�3a���������3j����$�6����$3��L�Lٌ�@z߰ߞ������5Pl�	P�A"//��;� e�P��t������P��O����w� ��S�>�w�b���B�/ ��������:(�J
�HZ    X��{�������2 E��� Ez��En.FZ���B��0,�1�0C��@�0� �?z���������/!/3/E/W/��DFp!����sq�����1�1�
  ^/�/�/�/�/	??-? ??Q?c?u?�?�?�?����5��fXst���K����1 @D���@�0?G�A � `?�AG�Ɛ�4�1<���;�	lB�}�RKLC@iK��F���2O�?�O����O�L��$H�O�O �$__H_3_l_W]�0�`@�_�W��_!��A���_�Xa_o]U+UyUoo=���To�fk c�Gтo�fb&�f�o�m�2�	�o}^u0  '� vo 2]_V��GҡOyAx�BU��| @e�t4C�F�B �
�C�.�,b7�m�.{�  �7�:�"�a�q� �B>���ÏU� �����=�87�!�/�>ua�0A`4�y�k��I�>L��T=�Au+���׏e)�G��3B�p?fff?�p?&�9�*� 6�G�	�D4�Ed�H ���HD�����ܯǯ  ��$��H�Z�E�~� ��g�����ؿO�q�s� ѿ2�ͿV�A�z�eϞ� �ϛ��Ͽ������� @�+��_s�9ߚ����� ���U���*�<�۟ Q�c��ߖ������
��T��iX� ��;�&�ϕ�o%���q� ������������( L7p�m�� �����H 3lW�{��� ��/�2//V/A/ z/e/w/�/�/�/�/�/ �/??@?R?=?v?a? �?�?�?�?�?�?�?O O<O'O`OKO�OoO�O �O�O�O�O_�O&__ J_5_G_�_k_�_�_�_ �_�_�_o"ooFo1o joUo�oyo�o�o�o�o �o�o0T?x@�u����w(�q������&� �J�8�n�\�~����� ȏ���ڏ���4�"�J]�P̒Pf���b� ����x��ş���ԟ ���1��U�@�R��� v�����ӯ������`� *���3�5�G�}�k��� ��ſ���׿����pC�1�g�u�  2� �ϭϿ���������+�=�K���o߁ߓ���߷��������
 ����D�:�L�^�p� ����������� ���b����{J��_�+�[�H� �@D�  \�?�>b� � `?��h����C]�\�X��� ;��	lh�c�}�����l�����F��a�����+���� .�Є�N	�߄o ����]�����0]�Y�.�@N8�r�+UUwz=��ʹ�`�0X���a&f/-�N�[�:/�u0  '`/n(a�/��/`�u��/�(B �/> @� 45�!ECw��/[?�/?j?��?�?��0�?�7 � ȗ2:�S��!�%h��<O#O�?C .�YOkK�18�0�O�J>�I�p�:�?�O�/)�>L�Sĝ0A��ODO�O<O�3h��N�h�10?fff?40?&nP�?�_�4 u�iQu��9d��_b��_ SV��_oo<o'o`o Ko�ooo�o�o�o�o�o �o�o8�_�_�_1 �-������ �4��X�C�|�g��� ��%ӏ����U�y B���f�x�����;_�� ß]������>�)�[A0A�f��n� w�6�����/U7/��� ѯ
����@�+�d�O� ��s�����п�Ϳ� �*��N�9�r�]�o� �ϓ��Ϸ�������� 8�J�5�n�Yߒ�}߶� �����������4�� X�C�|�g������ �������	�B�-�?� x�c������������� >)bM� q������ (L7p�m� �����/�/ H/3/l/W/�/{/�/�/��/�/�/?�/2?7($1���T?f;P? �?t?�?�?�?�?�?�? �?(OOLO:OpO^O�O��L��P,RP�N Q ¤%?�OI8�O%__I_ 4_m_X_�_|_�_�_�_ �_�_o�_3ooWo�O ���o䈓o�o�o�o�o �o%I7Y�m����w  2 Ro���1�C�U�g�y��������ϏᏀ���)�HoM�[�
 [�:��O������ П�����*�<�N��`�r��B{���{JM�������B��� @D�  ��?}�£ � `??��Ȣ?�C�����F� �;�	lȢ�A}����̠)�E�F�ê��6���A�� |���E�䨮�i�G�� Ͽ��,�ͽ� �Q�`_ǽϹv��Р�p��!����+UU����=����&���`6и�@�N���&fd��vݮ��y��=�u0  '������������բa�9��B <W�� @����EC�A��������������-�;�  ���:o��qU�	�uȢ��q����� �@������8������>5ѩ�С��09�+S>L>ѳt��A�D��B�����Ȣ��Ȣ��?fff?��?&� ��� ��բ�դ��ĥ$¨ D���xc�� ����///>/ P/'/t/_/�/13 �/�/�/??:?%?^? I?[?�??�?�?�?�?  O�?��3O�?ZO�/{O �/�OO�O�O�O�O� _#_�OV_A_z_e_�_��_Am�A��T� �S�_�_�_�Z����_ Fo1ojoUogo�o�o�o �o�o�o�o0B- fQ�u���� ���,��P�;�t� _�������Ώ���ݏ ��:�%�7�p�[��� �����ܟǟ ���� 6�!�Z�E�~�i����� ��دï��� ��D� /�h�z�e�����¿�� �ѿ
����@�+�d� Oψ�sϬϗ������� ���*��N�9�r�]� oߨߓ��߷������ ��8�J�5�n�Y��}�=(��������� ������
���.��>� @�R���v���������(����eP�P&=A"d��V��[�p ������  K6oZ�~� ^ O�DH��/=/ +/a/O/�/s/�/�/�/��/�/?�/'?7  2�[?m??�?�?�? �?�?�?�?JJ?/O AOSOeOwO�O��O�J
 �O�G�O_ _0_B_T_f_x_�_�_�_�_�_"�O��{�J��$PARA�M_MENU ?��U� � DEF�PULSE�[	�WAITTMOU�T/kRCVBo �SHELL_�WRK.$CUR�_STYL-`�nlOPTA9a�oT�B�o�bCioR_DECSN:`�l�o �o1,>Pyt ������	�a�SSREL_ID�  �E1��U�SE_PROG �%j%�j��C�CRF`*�1c}�_HOST !j#!����w�T7 ���ۃ����݃�v�_�TIMEDb*���~`GDEBUG(��k�GINP_F�LMSK@�o�TRv~� q�PGA��5 _��I ����CH}�  q�TWYPEl@� �4�]�X�j�|����� ��į�����5�0� B�T�}�x�����ſ�� ҿ����,�U�P� b�tϝϘϪϼ���q�WORD ?		FOLG-c�	U�	MA�KRO+�SUCH�L�C2�S7T�T�RACECTL �1��Ua
 ��@� ��@ /s t{�2����ߩ�S�DT Q���U��o�D �� 	�1	u��ԋ�ԗ I��E��Ԏ��B���M��@�`��6���7 �И��!��Q�ҝ���S��F`���U��V��W��X��ҏ�ԏI��ԕ�I�Z�Җ�ԖI䖫 �Ґ��\�ғ��ԑ��_��`��a���b��c�Ғ�Ԍ4�J���a��/��J�/�*�z�.��.��+�+�s�-�
+��+�+�+�+��+�*�-�+�+��+�+�+�+��+�+�+�+��+��@-�+�+��+�ސ-�!+�"+�#�+�$+�%+�&+�'�+�(+�)+�*+�+�+�,+�-+�.+�/�J�
�ӧ J�  �� �R� Z� b�� j� 	�r� z� � �� �� ���R� �Z��b��j��� �r��z������������g��g ��g��g��gg�
gz1�z9�z�)�zI�zQ�zY�z�a�zi�z��	U��ԔI�@��@I���	A��B!&J���0��������	F��
�������"	G*��GI�H��HI�2�	I��II�I��J���B	K��R	L2��M��b	N��r0��z�Ђ	O�֒\�К� 0��1��UP��PI�Q��TI6�J�f�ԁ��6��7��҂�ԃ��9�҄��ԄI�;��<�҅���=�҆�ԆI�?���@�Ԙ`�Ї�ԇ
I��ԈI��`��'���Щ���� ׮+� �/D�/Dڪ/D�/D�/D�/Dު/D�/D�/D�/D�/D�/D�/D�/D�/D�/D�/D�/D�/D�+�Y�a�i�&1�&9�&)�&�I�&Q�&Y�&a�&T�F�&q�&y�&��U&��&����q�U�y���	��4�P:�)�T!�4�4 D�Ԙ�PJ����V:�)��I��Q��Y���a�1� � e>4�#`�0m o��#`J�#`��#`J� #`R�#`Z�#`b�#`j� #`�#`r�#`z�#`�� #`��#`��#`��#`��#`��+cZa�0�b:�d�0�b8�dz0�br0�b5�d:#`�!�a2�d� �bb �bZ �b R �bJ �b� �b"#` *�a* �bb �b���b ���b���b���b���bH���b��f+@�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�/DU�/D�/D�/D�#E �uo���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ ��uk����� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?OO+O=OOOaO sO�O�O�O�O�O�O�O __'_9_K_]_o_�_ �_�_�_�_�_�_�_o #o5oGoYoko}o�o�o �o�o�o��o1 CUgy���� ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i�{������� ÿտ�����/�A� S�e�wωϛϭϿ��� �������o=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� ����������1 CUgy���� ���	-?Q cu������ �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?1�?�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y�����s?�� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� ��'9K]o� ������� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o ��1oWoio{o�o�o�o �o�o�o�o/A Sew����� ����+�=�O�a� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q��c�u��$PGTR�ACELEN  �v�  ���A`ȋ�_U�P �����������y����_�CFG ������Aa����� �ĝ�����������DEFSPD e���@a��Ћ��IN��TRL ɟ����8��V�PE�_CONFI���>�������]#�LID�á�����GRP 1���� ��v�C�  ��f�fAaA�\)G��ŎG�G��tA�  D	-��zA`d��)��9��� 	 �����S� ´  B��n�ے�������������B'?]�B�%��G��Y�C� <t�<��^���Z����� ������v� 9��I�oZ�%�����
� CDۿ���@� vA��=I~�H�?�HI;���� ��=(Ms�^ ���<���z�v���/�^�!��
V7.1�0beta1�� @j�H@'?�@,����B!�C�  C�\ .�T#D��k!_T#E�0` E) D�`g CH ��C/\ ~��C�� Ap�����BPffC߰ffAް ٙ�B(ffB<� A �#B<� ��33������? �§4����/?���&�8�����[?�?j?�? �?�?�?�?�?�?!OO EO0OiOTOyO�O�O�O �O�O�O_�O/__,_ e_P_�_ܳ �_�_n_ �_�_�_oo=o(oao Lo�opo�o�o�o�o�o��./T#F@ `>y:}N`|~ ?� �&������/�? ?/?A?J��on���k� ����ȏ���׏��� �F�1�j�U���y��� ��֟�ӟ���0�� T�?�x����_����o� �ϯ��,��)�b� M���q�����ο��� �1c=�O�y� ��ϸ������	�� -�?�H��l�Wߐ�{� ���߱��������2� �V�h�S��w��� ���������.��R� =�v�������[����� ����*N9r �o����� �/�a�;Mn�ϒ������$PLI�D_KNOW_M�  :%��>!�SV ����������)/;/M/�@q/\/n/�/�� ��M_GRP 1�\�� lC��"�$�`	`l�& �z0[��@�( "1*5&?8<���	7�+ a????�?S?e?�?�? �?	O�?�?9O�?OuO�+D�MR�#��-T���� ��O�N _�O�O6_�O
__._ �_j_d_v_�_�_���{ST�!1 1���"`� 0V�aciarC.�����@�y�pAßnIn��H���I,��sCon R�ep. Pies�:c7<j��F�@��gA�k�I��H��
�I0�]b.�P. y Dia�. an`� ���a�@��NA��*�IO�H���I1i�Llen1lD�����@� v�A�=I~��H��HI;��s]a�`dem1e�C/  �D��@��A����I�H���_I,���� �" 3�-?Q�u@���� o�!2o)`� �C��8�J� x�n�����ӏ��ȏڏ ����"�c�F�X�j�@���������k3� (��̟-�n�Q�c��� ������������4� �)�;�M���q���Ŀ������c4�'�� ˿,�m�P�bϣφϘ� �ϼ�������3��(� :�Lߍ�p߂��ߦ߸ߔ��c5�&���<)�n6�%�7�I�c7b�t���c�8��������cMA�D  �$"c � dPARNU�M  ��"|��7�T_SCHN� \�
��o�����UPDo����!>b_CMP_� Q����'�S_E�R_CHK6����cO3ERS8�@��"_MOP���_��RES_�G`�� ?aD^�-�B�}�Iw�(A.���oaDf��(B�I�8�4�1�V � Dh�RiHB�7Iw��9T2� ��`D�-?hC���I���t>�h  pD]����B��I��K�.�+ 2�VK ����/�//�	 ��1//�/y/�/�/ �/�/�/?�/(??L? ??Q?p?6/��Q/�? u?�?�?	O�?-O O2O cOVO�OzO�O�O�O�O �?���?�O�OD_7_ h_[_�__�_�_�_�_ �_
o�_o.o�O��\_Qo�a�no�o �o���o�o�o�����o�V 1���������^��`�^h�]��T�]���THR_INR� S���d�d�vMASS6� Z�wMN��s�MON_QUEU�E �š�����%MJ� 2���y��4A� 3 @��Bʡ��	�N- UqN8�v_m�ENDo�����EXE������B�E��y�j�OPTI�Ov��m�PROG�RAM %�z%�l�J3�k�TAS�K_IP�ߎOCFG ���󔟛��ODATA�1��}�@��"Ғ2/ ޖ�ߗ��
)�	����	������ې EF�<P�G�G�f��G�P�7N�= -� / 0 ; %? D F G1�4���J����ǭ����Y���m��ڑ3	��&�0�B�X*�T�>�B�G����&��������ϱi� C������������d�B�b���n� ��ҿ������ڿ6�*� F�`�\�F�XϪϲߦ� �߲�����8�4�߀n�Lߊ�z���s�I�NFO���}����
��.�@�R� d�v������������� ��*<N`r*��I���� _@f�s���DIT ��}�@mU����WER�FL��rs��RGA�DJ �}�A�  '?��3�q�m�x��U��?C�ё<@�����%qq���I�dJ��U˒���\9fqrbbA�<t�t$&*z /" **:""���/'#UL"G%��!Q)Q���q/ sE/W/i/{/�/�/�/ �/�//?�/??�?�? S?e?w?�?�?�?�?�? �?�?OO+OUOOOaO sO�O�O�O�O�O�O�O __'_9_K_]_�_�_ �_�_�_$o�_�_�_o ko5oGoYo�o�o�o�o �o �o�o�o;1 CUg����� ���	��-�?�Q�`c�u������ 	�� ,��P�;�	)u�#A� ��=�Ɵ���
// �@/ʏ܏q� ���L� ^�˯���������ܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�Dϱ�h�zό� �����������N�� .�@߭�d�v߈ߚ�� ����������*�<� N�`�r������� ������&�8�J�\� n�������������G ��"4�Xj| ����
C.l� v<�8�؟��� � �2������ >/P/b/t/�/�/�/�/ �/;?�/??(?~?L? ^?p?�?�?�?�?�?7O �? OO$ONOHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_o�_�_�_
owo .o@oRodo�o�o�o�o �o�o�os*< N`������ ����&�8�J�\� n��������#��G� ^h����R���ş� � /*/�6/��ҏg� ����B�T�~�x����� ����ү�����,� >�P�b�t��������� ο�M���(�:ϧ� ^�pςϔ��ϸ����� I� ��$�6ߣ�Z�l� ~ߐߺߴ��������� � �2�D�V�h�z�� �����������
�� ��@�R�d�v������� ����&���< N`r����  9Kb�l���.����$PRGNS�_PREF ����� �� 
�IORIT�Y  ݔ�����MPDS?PON  ݖ���#UT&�5&�ODUCT_ID' �"���OGGRP_TG�L$m&V&TOEN�T 1�i*�(!AF_INEE ��/�!tcp|�/�!ud�/~�!icm!?��Z"XY_CF�G ��+ ��)� #��?�?� ��?�?�5�?�?�? !OOOWO>O{ObO�O@�O�O�O�O�O_*Y#t3�� %�O_a_^�>�%a�#�!/�:_�_��-%�X��A���,  ���_
oo.o)(�T����0"�PORT_NUM#�� %�_C?ARTREP& {<��SKSTAE' ��jSAVE ��i*	2600/H620���!�_'3?K 	�ox����ݓe@������
�|�JU��e_�  1��+ p��������"�������a__CONFIw0�Zg #�]�U�ޔ��0蒯���ȃPt22�֋���[��C�U��$L�q�2�։�a����W8���p���k��?b?��̿XFN9D�v?W�g?�� =�2D����D4��D���������ɟ)#ݑ?��V�p�� B�4��ݑ� y���i�����_���� ��_��U]��A���Q� w��ۯ�����#��� �Y��=�˿)�sυ� ׿鿻�������U� ��9�Kߝϯρߓ��� �����������c߭� G�Y��}���ߛ��� ��)�s�����C�U���y�����k2S_M�OTI$ 2�֋
��=l�a0!@{�	��RUP90Y3?��%$��.#^,0047�K� =~�Y	�	������� D�~�D]�D!�^/����� d��i���D^L)D"��ݑ>>�?�b����|�?�^�=ڲO>���+>�c���%�@�	��O����LDw(U�J!�^A�`��Z  �����T����� �dstt 
+=Oas� �����a9���޵��x�	t �� /2/D/V/h/z/�/ �/�/�/�/�/�/6����3Dd?=?O?a? s?�?�?�?�?�?�?�? OO?"?KO]OoO�O �O�O�O�O�O�O�O_ #_O0OBOk_}_�_�_ �_�_�_�_�_oo1o Co>_P_yo�o�o�o�o �o�o�o	-?Q Lo^opo����� ���)�;�M�_�q� l~����ˏݏ�� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ��կ�����/�A� S�e�w����������� ̯����+�=�O�a� sυϗϩϻ���ȿڿ ���'�9�K�]�o߁� �ߥ߷����������� #�5�G�Y�k�}��� �������������� C�U�g�y��������� ������	�(�Q cu������ �)$6Hq �������/ /%/7/I/DV/�/ �/�/�/�/�/�/?!? 3?E?W?i?d/v/�?�? �?�?�?�?OO/OAO SOeOwOr?�?�O�O�O �O�O__+_=_O_a_ s_�_�_�O�O�_�_�_ oo'o9oKo]ooo�o��o�o�i�Q�d�P ��d@o���Q%?UP903�h�o��b$�b.u00+40�bQ�P�d�b�	�	��Q�a�b� D��D]��.D!���˨��Pd�RYr���D^L)D"��8�>CP�?b�B��y��?^�=ڣ%�>���>�b����#׿@����O�X��j�D$
�Q�^I�<y�R�P͟ 
 �a�P�����Q �dstt �o	��-�?�Q�c�u����������Ϗ�h�s.�v�sX�y�� 0�B�T�f�x������� ��ҟ䟟_�_�_,�>� P�b�t���������ί ������:�L�^� p���������ʿܿ�  ����1�Z�l�~� �Ϣϴ����������  �2�-�?�h�zߌߞ� ����������
��.� @�;�M�_߈���� ��������*�<�N� `�[�m���������� ��&8J\n �{�������� "4FXj|� ������// 0/B/T/f/x/�/�/�/ ���/�/??,?>? P?b?t?�?�?�?�?�/ �/�/OO(O:OLO^O pO�O�O�O�O�O�O�? �?_$_6_H_Z_l_~_ �_�_�_�_�_�_�O�O 	_2oDoVohozo�o�o �o�o�o�o�o
oo @Rdv���� �����%7 `�r���������̏ޏ ����&�8�3�E�n� ��������ȟڟ��� �"�4�F�X�S�e��� ����į֯����� 0�B�T�f�a�s����� ��ҿ�����,�>� P�b�tφρ������� ������(�:�L�^߀p߂ߔߢڬ��԰� �����?3T��@�f.%U�P903���߬�%�$��.��004�1��T���Դ�	��	���@v�`�����D�yD�^�CD!̴����V��d��I�����D^L)D"��8�>�@z?b����w^?^ =���>���>��c �� �@����P��?Z�D!��������ѯ�  �
��  ��љ������dsu
 t������/� A�S�e�w���������ʪ���
����w~�� ds�� �� 2DVhz ������ϡϳ� .@Rdv�� ������*/ </N/`/r/�/�/�/�/ �/�/�/?�/!/J? \?n?�?�?�?�?�?�? �?�?O"O?/?XOjO |O�O�O�O�O�O�O�O __0_+O=OOOx_�_ �_�_�_�_�_�_oo ,o>oPoK_]_�o�o�o �o�o�o�o(: L^pko}o��� �� ��$�6�H�Z� l�~�y���Ə؏� ��� �2�D�V�h�z� ��������ԟ���
� �.�@�R�d�v����� ������˟����*� <�N�`�r��������� ̿ǯٯ��&�8�J� \�nπϒϤ϶����� տ���"�4�F�X�j� |ߎߠ߲��������� ���0�B�T�f�x�� ������������� �'�P�b�t������� ��������(#� 5�^p����� �� $6HC U~������ �/ /2/D/V/Qc �/�/�/�/�/�/�/
? ?.?@?R?d?v?q/�/ �?�?�?�?�?OO*O <ONO`OrO�O�J�1�D��0 �D@�7��1%UP90Q3�H�O�B$�B.�O^�E0042�BY�0y �D�B	�	��1��A�B D���D^6.D"A_"�����0d�2�9R��D^L)D�"�8�>�4?b�����v�?^�=�ک�>��6>��^�����@���Q���&D-�1τ^?`Y�0 ��0�  ��A�0-�0��1d2 t�O�_�_oo /oAoSoeowo�o�o�o��J�P
 �W��Ġ1 ds �P�_�o"4FX j|����?�? �?��0�B�T�f�x� ��������ҏ��� �,�>�P�b�t����� ����Ο������� :�L�^�p��������� ʯܯ� ����H� Z�l�~�������ƿؿ ���� ��-�?�h� zόϞϰ��������� 
��.�@�;�M�v߈� �߬߾��������� *�<�N�`�[�mߖ�� ����������&�8� J�\�n�i�{������ ������"4FX j|�������� �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/���/??(? :?L?^?p?�?�?�?�? �?�/�/�/O$O6OHO ZOlO~O�O�O�O�O�O �O�?�? _2_D_V_h_ z_�_�_�_�_�_�_�_ �O__@oRodovo�o �o�o�o�o�o�o o%oN`r��� ������&�8� 3En���������ȏ ڏ����"�4�F�A� S�|�������ğ֟� ����0�B�T�f�a� s�������ү���� �,�>�P�b�t����������%UPg022��ɿ%$��y.��0013���!ʽ	�
Τ� ' �������)��D�D^L)�D"�8��>?V�G6j��v���<����,�p�׌��&�?65�������(�?�ø��C�>h����^=씵8�� ����� ������d2���������� ��1�C�U�g�yߋߔ�߈���
����� dst������%�7�I� [�m�����p��� �����!�3�E�W�i� {��������������� /ASew� ��������� +=Oas��� ����/�9/ K/]/o/�/�/�/�/�/ �/�/�/?//0/Y? k?}?�?�?�?�?�?�? �?OO1O,?>?gOyO �O�O�O�O�O�O�O	_ _-_?_Q_LO^O�_�_ �_�_�_�_�_oo)o ;oMo_oZ_l_�o�o�o �o�o�o%7I [mzo�o��� ���!�3�E�W�i� {�������Տ��� ��/�A�S�e�w��� ������������� +�=�O�a�s������� ����ȟڟ��'�9� K�]�o���������ɿ ۿ֯��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� ��?�Q�c�u��� �����������)� $�6�_�q��������� ������%72� D�m����� ��!3EWR d������� ////A/S/e/r)||r�%�)%�&�/�)��/�/�/�%p�% � �/?r8�?U?g?y?� l~�?�?�?�?�? O#O5OGOYOkO}O�O b�?�O�O�O�O__ 1_C_U_g_y_�_�_�_ �O�O�_�_	oo-o?o Qocouo�o�o�o�o�_ �_�o);M_ q�������o �o�%�7�I�[�m�� ������Ǐُ��� 
�3�E�W�i�{����� ��ß՟������ A�S�e�w��������� ѯ������&�8� a�s���������Ϳ߿ ���'�9�4�F�o� �ϓϥϷ��������� �#�5�G�Y�T�fϏ� �߳����������� 1�C�U�g�b�tߝ�� ��������	��-�?� Q�c�u��������� ����);M_ q��������� %7I[m �������/ !/3/E/W/i/{/�/�/ �/�/���??/? A?S?e?w?�?�?�?�? �?�?�/�/O+O=OOO aOsO�O�O�O�O�O�O �O�?�?O9_K_]_o_ �_�_�_�_�_�_�_�_ o__GoYoko}o�o �o�o�o�o�o�o 1,o>ogy��� ����	��-�?� :Lu���������Ϗ ����)�;�M�_� j�l�b�x���%s����� ��͟������<`���  ��b�8�E�W�i�� \�n��� ��˯ݯ���%�7� I�[�m��R�����ǿ ٿ����!�3�E�W� i�{ύϟϚ������� ����/�A�S�e�w� �ߛ߭ߨϺϺ���� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ����������#5G Yk}����� ����1CUg y������� 	/(Q/c/u/�/ �/�/�/�/�/�/?? )?$/6/_?q?�?�?�? �?�?�?�?OO%O7O IOD?V?O�O�O�O�O �O�O�O_!_3_E_W_ ROdO�_�_�_�_�_�_ �_oo/oAoSoeowo r_�_�o�o�o�o�o +=Oas��o �o������'� 9�K�]�o�������� �ۏ����#�5�G� Y�k�}����������� ҏ����1�C�U�g� y���������ӯΟ�� 	��-�?�Q�c�u��� ������Ͽ�ܯ� � )�;�M�_�qσϕϧ� ������������7� I�[�m�ߑߣߵ��� �������!��.�W� i�{���������� ����/�*�<�e�w� �������������� +=OZ�\�R�h�t	%c��HI��  stP�t  ��R�8�5GY� L�^��� ����//'/9/ K/]/o/B�|�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�/�/�?�?�? �?OO1OCOUOgOyO �O�O�?�?�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�O�O�_oo)o ;oMo_oqo�o�o�o�o �o�_�_�_%7I [m����� ��o�o!�3�E�W�i� {�������ÏՏ��� ���A�S�e�w��� ������џ����� �&�O�a�s������� ��ͯ߯���'�9� 4�F�o���������ɿ ۿ����#�5�G�B� T�}Ϗϡϳ������� ����1�C�U�g�b� tϝ߯���������	� �-�?�Q�c�u�p߂� �����������)� ;�M�_�q�������� ������%7I [m�������� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/���? +?=?O?a?s?�?�?�? �?�?�?�?�/�/'O9O KO]OoO�O�O�O�O�O �O�O�O_OOG_Y_ k_}_�_�_�_�_�_�_ �_oo_,_Uogoyo �o�o�o�o�o�o�o	 -?JcLaBaXudy1%Sv}�w t���qd}ds@cdu  q��Ba8��%�7�I��  <oNo��������Ϗ� ���)�;�M�_�2o l�������˟ݟ�� �%�7�I�[�m��z� ����ǯٯ����!� 3�E�W�i�{������� ��տ�����/�A� S�e�wωϛϭϨ��� ������+�=�O�a� s߅ߗߩ߻߶����� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� �������������1 CUgy���� ���	?Q cu������ �//)/$6_/q/ �/�/�/�/�/�/�/? ?%?7?2/D/m??�? �?�?�?�?�?�?O!O 3OEOWOR?d?�O�O�O �O�O�O�O__/_A_ S_e_`OrOr_�_�_�_ �_�_oo+o=oOoao so�o�_�_�o�o�o�o '9K]o� ��o�o�o���� #�5�G�Y�k�}����� ���������1� C�U�g�y��������� ��Ώ��	��-�?�Q� c�u���������ϯ� ܟ��)�;�M�_�q� ��������˿ݿ�� ���7�I�[�m�ϑ� �ϵ����������
� �E�W�i�{ߍߟ߱� ����������/�:�<�2�H�T�%C�m�w����d�� 3�4T�T�0�T�  q����2�8����'�9��  ,�>�w����������� ����+=O"� \�������� '9K]oj |������/ #/5/G/Y/k/}/x� �/�/�/�/�/??1? C?U?g?y?�?�?�/�/ �?�?�?	OO-O?OQO cOuO�O�O�O�?�?�? �O__)_;_M___q_ �_�_�_�_�_�O�Oo o%o7oIo[omoo�o �o�o�o�o�_�_�_! 3EWi{��� �����o/�A� S�e�w���������я ������&�O�a� s���������͟ߟ� ��'�"�4�]�o��� ������ɯۯ���� #�5�G�B�T�}����� ��ſ׿�����1� C�U�P�b�bϝϯ��� ������	��-�?�Q� c�u�pςϫ߽����� ����)�;�M�_�q� ��~ߐߢ�������� �%�7�I�[�m���� �����������! 3EWi{��� �������/A Sew����� ��//+/=/O/a/ s/�/�/�/�/�/�/�/ ��'?9?K?]?o?�? �?�?�?�?�?�?�?�/ ?5OGOYOkO}O�O�O��O�O�O�O�O__����$PURGE�_ENBL  |,A-A�-A�4PWF<PDO  �DT,BOQ TR_I�]TgQKUTQRU�P_DELAY ��"A"AKU,B�R_?HOT %�UiR�%+B�_�]�SNORMAL�XKR�_!o�WSEMI o&oeopQ�QSKIP_GRoP 1ĞUMQ x 	 ho �o�o�o�o�o�i�U 'wGYk1�} �������1� C�U��e���y����� ӏ������-�?�Q� �u�c���������͟����)�;��U�$RBTIF^T�ZY�CVTMOUT^V��U�Y�DCR��cƈi ���a?�7� uB��OoDvd'B��|d�m��P��BpňCX ��o���;��;���y0���$;�UU;���p/@�j�{� {� ����ſ׿����� 1�C�U�g�����vϯ� �Ͽ�����	�L�-�?� ��c�u߇ߙ߽߫��� ������)�;���_� J��n������ � ��V�7�I�[�m�� ���������������� ��3WB{f� �����*�/ ASew������,kRDIO_T�YPE  �[���REFPOS�1 1Ǟ[
 x	SoY)�}/��/ �-L/^/�/�/�/?�/ A?�/e? ?b?�?6?�? Z?�?~?OO�?�? O aOLO�O O�ODO�OhO �O_�O'_�OK_�Oo_ �__._h_�_�_�_�_ o�_5o�_2okoo�o�*o�oNo�o�o/%2 1�;+J/�o�oL �opvo�/��� ����6��Z�l�-'3 1�
�� V�ԏ��������@� ۏ=�v����5���Y�x�p�0$4 1ʍ� ����۟Y�D�}����� <�ů`�¯��������C�ޯg���0$5 1���&�`�޿ɿ� �&���J��Gπ�π��?���c���z�0$6 1�;+�������`��τ��3!7 1��.�@�z������>��S8 1α��������x��/�SM�ASK 1�� pH ������XNO����4�D�/!MO�TE  �M�_CFG �[�D�."PL_RANGW��+!_���OWER �;%��g�."�SM_DRYPR/G %;*%X� ���TART ����
UME_PR�O����j,$_EX�EC_ENB  y�c�GSPDC ̅ �e��GT3DB��
RM��MT_��T��Y���OBOT_ISOLC����x'NAME ;*�KJBVTU�211150R0�1xB V#_O�RD_NUM ?���
!H�620  �89�5 	���jx� �/ �PC_TIMEO�UT�� x/ S2�32t�1�;%�� LTEAC�H PENDANP�p�G�I�nW����Mainte�nance CoGnso�C�R,"b/���	UnbenutztY*�/X/�/�/��/�/�/�b"NPO� �K���SoCH_LF ���	�1T;MAVGAIL��5��c��SPACE1 2=��
 K?H HG�v�F������~4L8�?�L; WOL?;O�O�O�O�O�G �?OO%O�OIOkO]_ ~_A_�O�_�Y�#��] �O__%_�_I_k_]o ~oAo�_�o�o�o�O�_ o!o�oEogoYz= �����o�o /�Suw9����� ��������+�ُ O�q�c����������� ߏ���'�՟K�m� _���3�������˯� ���#�ѯG�i�[�|� ?�������ǿ���� �1�C�U�WϾ�;ύ� �υ������	��-� ��Q�s�e�7߉ߪ߼��ߥ��52�?�?��� #���G�i�x��\�� ��������*�<�N� `�r�t���X������� ����&�8�J���n� ���T������ "4F�j�~ �R���� 0B�f�z/�/^/ ��/�/�///,/>/ �/b/�/v?�?Z?�?�? �?�???(?:?L?�? p?�?�?VO�O�O�O�O  OO$O6OHO�OlO�O �_�O�_�_�_�_�O_  _2_D_�_h_�_|o�o Po�_�o�o�o
oo.o @o�odo�ox�\������3��
� .@�d�����y� ˏ�ӏ�5�G�Y� k�}�������u�ǟ� �����1�C�U�g�� ������q�ï���ͯ �-�?�Q�c������ ����o����ٿ�)� ;�M�_�σ����ϸ� {�ݿ�����%�7�I� [�	�ϡϓߴ�w��� ������!�3�E�W�i� �߯߱�s������ ���/�A�S�e���� �������������� +�=�O�a������ �m����'9 K]����y ���/�4�'� 9K]/���/�/ �/�/	?�/?#R/d/ v/�/�/�/�??�?�? O�?O<?N?`?r?�? 2O�?�?�O�O�O__ �O8OJO\OnO�O._�O �O�__�_�_o�_$o F_X_j_|_*o�_�_�o �o�o�_�o BoTo foxo&�o�o��� ����>Pbt �4�������� ڏ�:�L�^�p���0� ��ȏ���ޟ����� 6�H�Z�l�~�,���ğ ��ׯ�������"�D� V�h�z�(�������ӿ@���	���#+52.D/V�h�z�(Ϟ��� ���ϳ��&��;�#+6O�a�sυϗ�E߻� �������"�C�*�X�#+7l�~ߐߢߴ�b� ����	�*���?�`�G�u�#+8������� ����&G
\}xd�#+G �5+� �:
�  �,:5% K]o��������o�>d �%/ 7/I/<j/|/�/�/� ���*�/�+?
/;? M?_?q?d/�?�?�?�/ �/�/�/?O7O*?[O mOO�O�?�O�O�O�?��?�?O$O6_ `� @> oU�}_ �O�_�Ek_9_�_-Oo �_�_�_�_loo1oSo �ogo�A�a�E�c�o�o !�e�oSe� 9k����������L
�_n�@�_MODE  �^��S ��]�_Z���_�9��	4�]�D�CWOR�K_AD�����F�R  ���b���_INT�VAL�������R_OPTION̖� ��F�TCFB� ۗ���?��7����V_DATA_?GRP 2��H�DU@PJ�y�F��� ��G�ʯ���ܯ� � 6�$�F�H�Z���~��� ��ؿƿ����2� � V�D�z�hϞόϮϰ� �������
�@�.�d� R�tߚ߈߾߬����� �����*�`�N�� r����������� &��J�8�n�\�~��� ������������4 "DjX��Be�� ������q�5# YG}k���� ���//C/1/O/ U/g/�/�/�/�/�/�/ 	?�/??-?c?Q?�? u?�?�?�?�?�?O�? )OOMO;OqO_O�O�O �O�O�O�O�O___ %_7_m_[_�__�_�_ �_�_�_�_�_3o!oWo Eo{oio�o�o�o�o� �o� ��o�oAw e������� ��=�+�a�O���s� ������ߏ͏��'� �3�9�K���o����� ɟ���۟�����G� 5�k�Y���}������� �ׯ���1��U�C� e�g�y�����ӿ���� ��	��Q�?�u�c� �χϽϫ�������� �o>�b�M�ߕ�� �ߧ���������� %�[�I��m���� ��������!��E�3� i�W�y�{��������� ����/eS �w������ �+O=sa ������// 9/'/I/K/]/�/�/�/ �/�/�/�/�/�/5?#?�Y?+��$SAF_�DO_PULS � -��������1t0CAN�_TIME�0}��3���1R �����8�	U	����
�8��U�4�4�� ^� OO0OBOTOfO�?�O��O�O�O�O�O�G]�1  B2TD�1�1dXQ Q�4q}��1�� @CV T[�0P_z_�\�1�_�W�P�U�� @=B�3T i_�_��_oiT D��oAoSoeowo�o�o �o�o�o�o�o+�=OaX^?VNV=py 
�qp��y�3�1;��o}��4p{}
�?t� �Di�0�A��1�z   �@B�1�q�1�A�1z��Y�k�}�������  �������� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����$��h_H� Z�l�~�������ƿؿ'�>T�Q���R� 7�I�[�m�ϑϣ���ρ�0�22�@U<�}����$�6�H�Z߁�^�^ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� ������������� ,>Pbt��� #�����(�:L�2��P��imih� �0�A�B Ѓ��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�?@OO*O<ONO#��=X ��*`YO�O�O�O�O�O �O__&_8_J_\_n_��_�_�_�_�Z�B�p�_�V�_i��A���_/m	123�45678�r`!B  �/h�@��jo|o�o�o �o�o�o�o�o q�O# 5GYk}��� ������1�C� T�w���������я �����+�=�O�a�ps�����V�BH�� П�����*�<�N� `�r���������̯ޯ<�[�:�j��&� 8�J�\�n��������� ȿڿ����"�4�F�]�D�_wωϛϭϿ� ��������+�=�O� a�s߅ߗ�Z������� ����'�9�K�]�o� ������������ �#�5�G�Y�k�}��� ������������ 1C�gy��� ����	-?@Qcu���Ug` ���`�//%(�"C��A�_J �  >%tA2qB�gb%)
�Pdq#�
?`��R2��/�/�/,�/�+pM$ZO���/0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O?�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_��_�_ ooG!�$S�CR_GRP 1����� �t �G!� R%	 _Ra�Zb kbdd�f%f!�ekwgp�o�o�o(-�a ��bD�@ D�@� =qcw�k<M�-900iA/3�50_iC 67�890� @t�a�M9A3NqC#
V06.10 zpD�h�a�br#�u�vZa�fIa�cIa3f!"�ahj�a�y	�r��
��.�@�P��G�H��r�r^g�v�P�0D�)��D�yzD��3��1/��~ǯ�Bd�vaA�������z���)@�7 @�*���K&P�  �=;��D�*5>��XD��Z`�OG!�o��o1�.'"��受hB�  B��|�z�����L ��  � q��va@���˟ ?���v�: 򟨛vaF@ F�`� %��I�4�m�X�}��� ��ǯ���n� q��h��m��4�B�E� گ��v�����ӿ��п 	���-��Q�<�u��/@���c�o����i
�����C#�@��"� ߘg�;� Z�R�?12345Or`��h���C$Aϐ�Ƴ�(㏛cd!2��G!A ��������2�>�P�� �v�(�|����  Ibp`�tZ`�}�{yi�� gϩo�iǑ�P������7uInde�pe��nt Axes Qs	����n �f�w��s�w3i� �r���j|��� �c��	�n�'9 ��Z��~��S� �w������/��� F/藦�t/��/��/ �/�/�/?�/?=?(? a?(�:�p?�?�?�9f� L?�?�?!OO1OWOBO {OfO�O�O�O�O�Or� ����`�A_��e_w_�_ �ONݺ_\�n�~�o ��L$o7o��boto�o Uo�o�o�o�o�o��S�����_� �:��._������� ��������p�$6 HZߏ���'�� ��o�~������Ho hퟀ��#��G�� h�
/��./P/R/d/� ��0�1��U�@�e� ��v�����ӿ�?�?� ����?Q�Ŀu�`ϙ� �ϽϨ��������� ;�&�_�
�_m��F_ X_�����_�_�_�_�V�_w�o����� �o�������+�=�� a�s���$6xBT ����3��W ���,�>�P�b�� ��������ΏSew ��:�L�^����/ /+/��ܟa/��/�/ 6��/Z��/~� ?��į ƯدZ?|/�?�/�?�? �?�?�?�?�?#OOGO 6� �VOhOzO@��O8O �O�O_�O1__A_g_ R_�_v_�_�_�_~�� �_L����Qocouo�2�8�J�8ff��o�� 4/Z�Wi8y����������$SEL_DEFAULT  �����P��MIPOWER�FL  6e.��7�WFDO#� �.��RVENT �1����,���`L!DUM_�EIP����j!AF_INE"�<Ə�T!FT��������!�>� ���e�!RPC�_MAINf�H��8T���x�VIS��G�y�����!TP�PU����d�I�!�
PMON_PR'OXYJ���e8�����c���f���!RDM_SRV�r��gЯ-�!RZ�dI���h�y�!
z��M����ih�ſ!?RLSYNCƿ��8���!RO�S��8��4 �]�!�
CE�MTCO�M^ϲ�kLϩ�!	�r�CONS�ϱ�l ����,�������B� g�.ߋ�R߯�v��ߚ� �߾�����?�����RVICE_KL� ?%�� (%�SVCPRG1�r���2����3������4
����5�2�7���6Z�_���7�������8������9������D������ '����O����w�� $����L����t�� �������?���� g�����=��� e���/��// ���W/��/��- �/��U�/��}�/�� �w������B?�? ��?�?�?�?�?�?�? OO?OQO<OuO`O�O �O�O�O�O�O�O__ ;_&___J_�_n_�_�_ �_�_�_o�_%ooIo 4o[oojo�o�o�o�o �o�o!E0i T�x�������M:_DEV ����MC:���n,%�~�L�   ���i��!�OUT�`�:�!�?REC 1�d5L���  M�� W	  �p �o �q �u�������㏔􍶃 �ۂ���ԏ5�D�
 �T�F�6��YU�h�	+�&M�FȀ�d5���� ��� ����M�#�� U� �97��7�Y7��~���,�� �  I7������ �DљUh_e6 ���3)����x�E�Yџ�K�K4�_ �-� 37��Z7��� v ��U�� �!j7� �	�����͐�}�V7���]����Ĳ�.�`��}� � � ���t��Vٯ > �7��7�j9�| ��� A ��k7�- �����u͐=���Q�	�����Gu��  ���$  ��}�)� ? ���=��X � �� d �QR7�� �7��͐����� ������u��u���չXGJEJa��.�K �e��$տ��� ��P ���P���7�W� �c7�����7�����1�� �27��7��7��}����FE��� ��� a ��M��� �YϪk�d7��7���� �<���M��͐�͐�j�}M����L!����P�
q��J �iM�z �t� ��H���V �sŴGj7�f �e��� ���͐��������Uܹ���J� ��߷�hM�� �* �/����ߔ�߾��M�͐@��UC�L7��U��ϰ��(� ��� �� Vl� �BQ�Y��P]�o�￢{吸j�������7�C���ca�	���rM�%��N��1��Z`���� �)��� 7��7���H�^R ������ H���������R�La�tp	��ZM�"�퐶}���%�u���� �|� � ����A �7�� ��7�� �:7��	��Q,9�j���� ��6�=�@
JѨ������	���4�*�M���S�E�M��M�2��?�^7�4  ����Z7����7����������� %��������� ��#5c����Ѥ��u�����dIO2<]�f��}�� #��  8�Ҥ�� @K4���E/ %g7�� � �7� ��.m/�������e�����ߋ���ڕ)M-�~
���}�$�e=}��N���4�/�O�5M�P�l �`ZM�S��\ �t7�f�� F7�,  j�/��� ��;� Mzj�A9R�X	�H��L�<  D�O��A?��H ��}�@� Un���? ȑ�7�U�7��7��7��?��xM���
���u����i:h4a	��j��P������V�? � �; ��y�������1�c�.������͐D�+��7�0�,:��XPP�ā�L�qOPё] �x������O��[-4�A(�,1����M�}͐�1���m�@��+}D��[
�S���}�J��kE_ ��R�����pO��T�7��L�_���� ����v]H��Q�c�u� ��������Ͽ�� .��o�o�o/SF���m�i��� ������!�3� i�W���{���Ï��� Տ�����/�e�G� u����������џ� ���=�+�a�O�q��� ���������߯�� 9�'�]�o�Q������� �����ۿ�#��G� 5�k�YϏ�}ϟ��ϧ� ��������C�1�g� y�[ߝߋ��߯����� ���q�Q�?�u�c� ������������� )��M�;�q���e��� ������������% 5[Im��� ����!1W E{]o���� ��////S/A/c/ e/w/�/�/�/�/�/? �/+??O?=?_?�?g? �?�?�?�?�?O�?'O 9OO]OKO�OoO�O�O �O�OI_E&__J_ 5_G_�_3��O�_�_�_ �_�_�_o1ooUoCo eo�oyo�o�o�o�o�o 	�o-Q?a� i������� )�;��_�M���q��� ����ݏ�����7� %�[�I����s����� ٟǟ����3��'� i�W���{�����կ� ɯ�����/�e�S� ����}������ѿ� ����O�_)�s�aϗ� �ϻϩ��������� %�K�9�o�]ߓߥ߇� �߷��������!�G� )�W�Y�k������ ��������C�1�S� U�g������������ ��	?Q3uc �������� )M;q_�� ������%// I/[/=//m/�/�/�/ �/�/A�k_$?g_H?3? l?W?|?�?U��/�?�? �?�?OOAOSO5OwO eO�O�O�O�O�O�O_ �O+__O_=_s_a_�_ �_�_�_�_�_o�_'o oKo]o?o�ooo�o�o �o�o�o�o�o# YG}k���� ������U�7� e���y�����ӏ���� 	��-��Q�?�a��� u��������ϟ�� )��M�?�?K����� ����ݯ˯����7� %�G�I�[������ǿ ���ٿ���3�!�C� i�Kύ�{ϝ��ϱ��� ������A�/�e�S� ��wߙ߿ߡ������� ��=�+�a�s�U�� ������������� %�K�9�o�]������� ����������!G 5kM_��������$SE�RV_RV 1�	8��0(	\��n���!3TOP10 1�=
 6 2q��g q��6��E sq� ��*"r _"$q�*�6 &q�F ��q�F *J!�YP�E  q���Hq�1HELL_CFG �8t&�0�? �?�/>q�%RSR�/�/ �/??:?%?^?I?�? m??�?�?�?�? O�?�$O5MDD<I�S �E%5OvO�OCE?Mbq��O�B�@�D�\D!d�Oq��)�}&HK 1�+ �O<_7_I_[_�_ _�_�_�_�_�_�_o o!o3o\oWoio{oC~}&OMM �/��o|"FTOV_E�NBi$Et*OW_?REG_UI�o{"�IMWAIT�b\�I{OUTvD�yTIMu���WVAL,s_U�NIT�c�vt%QL]CpTRYwt%�1MB_HDD�N 2�k �)P��bh��ICt{�����\\�ن�P��qۆI������[}h��E��N����8�q�<��7� I�v�m������̊�q�ON_ALIAS� ?e�iLhe p���(�:�L�D�� w�������X�џ��� ��ğ=�O�a�s��� 0�����ͯ߯񯜯� '�9�K���\������� ��b�ۿ����#�ο G�Y�k�}Ϗ�:ϳ��� �����Ϧ��1�C�U�  �yߋߝ߯���l��� ��	��-���Q�c�u� ���D��������� �)�;�M�_�
����� ������v���% 7��[m��N �����!3E Wi����� ��////A/�e/ w/�/�/F/�/�/�/�/ ?�/+?=?O?a?s?? �?�?�?�?�?�?OO 'O9OKO�?oO�O�O�O PO�O�O�O�O_�O5_ G_Y_k_}_(_�_�_�_ �_�_�_oo1oCo�_ Toyo�o�o�oZo�o�o �o	�o?Qcu �2������ �)�;�M��q����� ����d�ݏ���%��Ѓ�$SMON_�DEFPRO ����N�� *SY�STEM*Ѐ6B��>�RECALL� ?}N� ( �}׏����ԟ��� ���/�A�S�e� w�
�������ѯ��� ���+�=�O�a�s�� ������Ϳ߿񿄿� '�9�K�]�o�ϓϥ� �������π��#�5� G�Y�k��Ϗߡ߳��� ����|����1�C�U� g�y���������� ����-�?�Q�c�u� ��������������� );M_q� ������% 7I[m ��� ���~/!/3/E/ W/i/�z/�/�/�/�/ �/�/�/?/?A?S?e? w?
?�?�?�?�?�?�? �?O+O=OOOaOsOO �O�O�O�O�O�O�O_ '_9_K_]_o__�_�_ �_�_�_�_�_o#o5o GoYoko�_�o�o�o�o �o�o|o�o1CU gy����� ���-�?�Q�c�u� �������Ϗ�󏆏 �)�;�M�_�q���� ����˟ݟ��%� 7�I�[�m� ������� ǯٯ�~��!�3�E� W�i���z�����ÿտ ������/�A�S�e� w�
ϛϭϿ������� ���+�=�O�a�s����$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1z� �?��%�ߎ�������� @�G���E86�w���$f���0�������@�����s���7���%�f� �@� V���֐GX8�������������S����'���U�VY�$�� ؠ1����g����v���Sq}G�0�6w���f������ ל��8�/���1�7/�� /�&/g/�3q�e�/ ��R߆/��/�����/�/��c}��/'?�&����V?)�ACF?�?�קqv?�?�#7/�?�?�p�!�?O��E�OGO �X�86OwO�gyfO�O��?`�O�O���q?�O_�_O_�O7_�d��&_g_�GBy�V_�_JW����_ �蓰�_�_�1E�_&o �AaoVo� � Fo�o���n vo�o�c	�8�o�oւ���o��U`�Gjg�8�Ov �y�f���a5�� ���1���[G���7�����&�g���c�jV�����Eo�Ə�@��� �Y�1~�'��Gd��W��z��%��� ׆��v�����o��81;�_�����G�ƺw�6�w����8f����m20��ׯ�:?�Ư����1K��7�ֽ �f�� ד��V����w�q���ǿ�!(����֏�P�'��ǋQ��W� ���Fχ���1u���PA�RAM ����� �	�P�\�pb�������OF�T_KB_CFG�  ��ԉ�OP�IN_SIM  ����=�O�a�q`���RVQSTP_DSB&��߈�$SSR �)�� � & F�OLGE125 y.����0017a���Ī�THI_CH�ANGE1@�����GRPNUM�� �OP_ON_ERR��I�?PTN )���C�RI�NG_PR1�U���VDT+� 1�<����  	��* ����������0�B� T�f������������� ����,SPb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?k?h?z?�?�?�?�? �?�?�?
O1O.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\o�o�o�o �o�o�o�o�o�o" IFXj|��� ������0�B� T�f�x�������Տҏ �����,�>�P�b��t������VPRG�_COUNT�q�|��ƒENB�����M�4���UPD� 1���T  
����B�T�f����� ����ׯү����� ,�>�g�b�t������� ��ο�����?�:� L�^χςϔϦ����� ������$�6�_�Z� l�~ߧߢߴ������� ���7�2�D�V��z� ������������
� �.�W�R�d�v����� ����������/* <Nwr���� ��&OJ \n����������_CTRL_�NUMГ!��!"GUN%" 2�>0��  1$!�!f%#d'o/e&��/�/�/�/ÐYSDOEBUGА1�� �d�� SP_PA�SSЕB?;L�OG �0��� J1�^���k$[=�c%
M�C:\0413��12_7MPC6? 1$�)�]?o5UD1z52�.�3SAV �9=�!n- �8S�V�;TEM_TI�ME 1�R+ �( @�"0�n� "5v�,"hF�*sH@O�O�O�O�O�C�$T1�SVG S+�ѕ'���PASK_OPTIONА0��:ߑ'Q_DI0��ߔTBCCFG ��R+�=�.�_`�_���!�_�_�_ o�_5o oYoDo}oho �o�o�o�o�o�o�o 
C.@yd�������	��% �6��i�{��X��� ��Տ�����0��=P �!�G�5�k�Y���}� ����ßşן���1� �U�C�y�g������� ӯ������	�+�-� ?�u�[�F�������˿ ݿ[����7�%�[� m��Mϣϑ��ϵ��� �������E�3�i�W� ��{߱ߟ�������� ��/��S�A�c�e�w� ���������+� =���a�O�q������� ��������'K 9[]o���� ���!G5k Y�}����� /�1/��I/[/y/�/ �//�/�/�/�/�/? -????c?Q?�?u?�? �?�?�?�?O�?)OO MO;OqO_O�O�O�O�O �O�O�O__#_%_7_ m_[_�_G/�_�_�_�_ �_{_!oo1oWoEo{o �o�omo�o�o�o�o �o/eS�w �������+� �O�=�s�a������� ͏���_	��9�K� ]�ۏ��o�������۟ ���͟#��G�5�k� Y�{�}���ů���ׯ ���1��A�g�U��� y�����ӿ������ -��Q��i�{ϙϫ� ��;���������;� M�_�-߃�qߧߕ��� ��������%��I�7� m�[��������� �����3�!�C�E�W� ��{���g������� ��A/Qwe���� �$TBCS�G_GRP 2���� � � 
 ?�  ��� >(:t^��� ������/,/ /P/:/t/�/l/�/�/ �/�/�/?�/(?:?$? ^?D?n?�?~?�?�?�?��?�?O�?6OHMA���*SYSTEM�*� V8.230�6 qC4/2x@0�14 A t � _F_GF�� P�ARAM_T �  �$MC�_MAX_TRQ���$�D_MGNںCC� AV�IST�AL�IBRK�IN�OLD�FSHORTMO_LIM	Z��M�EJPTPL1�CU2CU3CU4CU5�CU6CU7CU8�A � �A��A�� �_ACCE�JR�WTQ�SPAT�H�W�Q�S�Q_RA�TIO�B�S�@ �2  	$CNT�_SCALE	ZS�CL�CIN�Q_U�CA��bCAT�_UM%hYC_I�D 	*cB`_�EKPGjTPGj]PG`P�AYLOAWJ2�L_UPR_ANG�fLW�k�a�i�a��ER_F2LSHRT�gLO�da�g�)c�g)cACRL_�Shpgzd�BHV�A`  $H��B:rFLEX7s�4�@Jb�@w :$aLENKQyguTQ$DEjx��t|s�R�X�p�zSL�OW_AXIqW$F1aI�s2�x�1�q�u�wMOVE�_TIMd_IN�ERTI%`:p	$�D	�TORQUEЧQ!��p�IHPACEMN�`��P�s�E^�V�p�A/�x�@�x�TCV���@��AP�������@T.�ሄ@��J�A����M�	�(a�(`J_MOqDa�p� R�*@�gq2�@P�^�!Eo�0`J��Xp�1A�RU�?�JK.���ڒ�KKSVKTSVK�]SJJ0�KSJJ�TSJJ]SAAKSA�ATSAA
�fSAAoS�AN1ǌ<����@��@PE_NUQ��VqCFG�A� � $GRO�UP�@SK&cB_CONFLIC�d�B_REQUIR�E.q�qBU sUP�DAT�v� �E�Lk� ͥ���$TJ�P�JE��@CTRa�qTN�	�F˦��HAND�_VB8rVqOPn�U $]�F2�F�
�TSCOMP_S�W&a�*Uq�F�� $$M�`�IR �C|��A��x��R���A_}b�FDļ�MA*�LA�LA�KA [Ұ��KD�LD�KD [Pf�PGR�Gp�ST�Ghp��Ip�NXDY�`R�@�E��ڵ�` `�g �q�g�a�g0�<Q@��p��UPKUTU]UfUoU�xU�U�R?�Vr�Tc r�Wt�R %�xn�TPy�ASYM�U:p� �V�Pm�ao_SHo�g4d]���C�>oPoboto�cJ��l>P�j^�T�i
�_�VI&���Ѫ�V_UNI�c��TS�aJ��������l���e ����m�y>P1�a���GtOs �(�TCPPIR�A�  ��ENAB�L�p����$TCDELAYݱ`����SPEE4P O X ��I�Nڠސ��ڠGP����Q����q�@MPڢPR�OG_���YPEtڡ��_z�	 |�m���SE s��m���|' ǦWARNI��sEN&���OTF�q�j��_T���MA�ARSCW����SPDz�
 ������?EARTBE��ѣET��z���PPAsRGAT��FLG�uT�|sS�@E�@R&�6�%�aos6�REAJVXTRx�OUT�A p렜��� E�̢F�ID`�(d^�Uc �A�`��޵�G�Qdu��PH���<�t�{I�$DO�� ���z�) ��I��A���J �p��W#�۠\���q�� � VT�MES���R�*��T P��"@P�l���#��(�!�)T�"�m� $DU�MMY1]Q$P�S_�pRF�pg@u$�&��FLA|���2�GLB_T`u�k*5����(����8!�����QSuTT��SBR�P�M21_V�T$_SV_ER�`O�Lp3�3CLD0p2A^�l���GL��EW�Ag 4��$��$ZݲW�3���`P�IAs %bYѵ1U�5� ]�N�0�w$GI�}$�1� ��1�0�A� L��F�}$FJ�EFN� M�NcyF]IJ�TANCb_  `�J RǱ� +!$JOI�NT�����3M$� �Q��FECE�q���S�bv*B���Q�� �pUS�?���LOCK_F�O�`[�� BGLV���GLXT  _X9M`�AEMP�@��� -PB2�@$US��!�0p2*��4QQ�RW��@QQ�SCE8j�CrP $K��}M#TPDRA�0�T�AVEClp�V�@kIUQQVQHE�@OTOOL�s�SV�t;RE�PIS3|s�T96*�)`ACH� ����QON��$29��"�PI�  @�$RAIL_BO�XE���ROB�O"T?�r1HOW�c>d� aROLM �"ge_�
dxb��/`�p�6�O_F��! !��0�Q^q�NY�R�PO]r�B�p�A"�`�A�2~X2MU��֡���@	 IP#VNK��R/b�Q
�QQ��`�PCORDED��@���`�A��OY  � D )0OB�٣�@dwSq�#E �Sr�ۡSYSSqAsDR =QTCH���  , �A��A_D�th�*�ޤAVWVA�� Ǥ �P�2kPR�EV_RT��$�EDIT�VSHWR����$�K��'IND� `;�$х�D&�[�U�6���KE��� �l�J�MPppLj/ RA�CE)[p�Ij,PSڢC �NE�P<ۡ��TICK�S���Mo�o ��HNR1 @]p��L	�_GK&f��STY�aLOD1_������~� t 

 G��u%$�qD=� SFp!$��8��!��F �P��LSQU�aLO���TE�RC� ݱZ�Sz� @h0�� p���㡼Q,�O� �#dI�Z4A��! Cx�"!�oUTPU���1�_DObB�pXS:�@KjAXIP��c�VQUR���0i#$ATH`�~vK���_�P�rET��P Rlp��%O�F��P�A������$ cc>  ���ĐR3� lѐu��A����� �������ù�ӹ R���R��R��d�~� B�d����҂�C翐��C��� �2�D�SY�ĐSC,0 ! �h�0DS�� X}�AT��<�� ~��~�"ADDRES�S=B�SHIF�HP�_2CH� zqI�K0���TXSCR�EEUr"	 k�T�INA�3@��Dp�񒡒�T0# T�� �0'�g00�^��r^�|�RROR_vA���(�h$�1UE5$$# ��Щq0S�1�q�RSM��T�UNEaX��j���S_�3���G�ѽ���G�C��B��� 1# 
z��%="�2��VMT!�Lv�m�rw0O�D�@UI_� }HP� & 8e�Bw@_T���f� R���Bcg�"� R�O���T0'���7$/BUTT��R Rra�LUM��u���ERV�R�Pa@��S1�({ ƠGEUR�&SF���A)� LP$���E��C�)#�S��1�c�1��P0�5.�6
.�7.�8�����a@���%�Q�ASv�'R�USR�4O) <Z0� UBr�AI΀@FOC�Q.@PRIΡm`��� TRIP�m��UN$ 5$*	@ t�$ kcjQ�IQ����� +a��� �G� \��1���\O	S�qR��V�H�QS1,�?�3�>���HRU�S1-����8��HOFF!PT0�.[p�O' �1,�09-�0G�UN_WIDTH|���B_SUB�"�p0�SRT� �/0��vA�` �OR`�'RAU��T�����VCC�М�0 ��aC36MFB5124 ��VC/0.D1h %bTq��A�4.��c)�C�`^	%DRIV���C_Vu�,$(��@D��?MY_UBY��$ V�vA�� B�tC�#�Q�tBi0pp+��"L7�B�M�1$��DEY�!�EXG�n��Q_MU��X�10orb����GðPACIN΁}�RGC�52�`2�32���!RE{����Q����2�0�2�TARG�@P�1Rc0��R� �03s d��_�FLA΀�r	�"N�RE�#SW0_A1 �@�!�O���A���3�EE��UB�a �`V�HKG�4���:`����05�!CEA��+GWOR!P�5���MRCV�5 ����OS�M!PC2S	phB`3hBREFF� �FqF\A�0�࿣�0�� mJ�A~J�A�K�EqFO�_RC,KXEKV�S����']#���6 �$���1؄��b%�pROU�[2�#O 1z52�2�Pa$���� �΀3��t2���Kq�SUL��c4;r��� 5�  �P@�3�cN�f��f��c�PL�#5e�#5e���Ag���$��7�0 &��ǡ4� 2��C�`+�LO�A�d@�a� �iu��`ܓC�p[MI��FR�hTj���fR[$HOh��r��`COMM'#��O�B�v{X���؇V�P]2�Hq_SZ3dcQu6/cQu12��`Nx0Lx�`LxWA�e�MP�zFAI�`G�T�`AD�y�!I�MRE~T�r_�G�P��� ��&ASY�NBUF�&VRTaD���qσOL��SD_�:�W�P�'ETU�#�`Q�0��ECCUP8VEM�:0�e���gVIRC��q2�T@#�8^P��0CKLAS^	��VLEX��9�/�����	�LmDLDE�FI<�� �r�������T�p�Q��:����T�1�'�����9V�� ;`��L����{,�"UR�3�0_R�p󔟑�!���U3 �/�/�$�`7���0Ғ� �TI�Q��SCO�� �Cz�4;#6; �;�;!�;/�/ /%*ᢕ���D�S�^�@ �_�M#<)���J*��%��q�=)G�egLIN���W�@sXSGAq�>  ���N�BPK�cH��HO�L�� ��ZABC}?v2`�XS��@
 ��ZMPCF}@<����ԙ��l!LNI�΀
q���� ~A ���xq+@��CMCM0}CKsCART_ٱ�#�P_�� $J���������pS��S��2UXW� ��UXE�!A�<��9��d�J�\�J�lƿ ��ZPץB� ��b"�h��Y:!�D" Ca⣖��IGH&3G�?(!�!��A� ���D � T��A~��$B�PK�'E@K_Xa�	c�RV�`F���Ba�OVCY��籠�TU�O0��j�
RI��1uD��TRAC�Ex�V
1���SP�HER��E ,�!�������|�$T�b� 2������ �dX,�?� �	 HD|�9 ��'�L��0�)�?D�fAp�M��Z�D��'�9���BHZ�\�n��\�����C���f�ff���CA�fB����������I�H3�����z���@� H�I����������&�C n��pP��	V3.00~�	m9a3�'	*� �����J�𙙚�x�dp	 �   @��]2f�x�� �� �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?O��	 O2O O^OlI0pO�ODlO �O�Kz�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>PbO >O�JO���O��O �(��O0�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯t ���.��B���v������J�� ���  Vf���2f������	 2?�*�c�Nχ�rϫ� �ϻ��������)�� M�8�q�\�nߧߒ��� ���������#�I�4�m�X��|������ ��������8�#�\� G���k����������� ����"XC| ���I�s���� �!E3UWi �������� /A///e/S/�/w/�/ �/�/�/�/?�/+?? O?a?k��p?�?�?>? �?�?�?�?�?OOBO 0OfOxO�O�OZO�O�O �O�O�O_,_>_�O
_ t_b_�_�_�_�_�_�_ �_oo:o(o^oLo�o po�o�o�o�o�o �o $H6X~l� ������?�&� �?�h�V���z����� ���ԏ
��.���� d�R���v�����П� �������*�`�N� ��r�����̯��ܯ� �&��J�8�n�\�~� ����ȿ���ڿ��� 4�"�D�j�Xώ��:� ����tϢ�����0�� T�B�x�fߜ߮����� ���������P�b� t��@�������� �����L�:�p�^� ��������������  6$ZHjl~ ������ 2 ��J\n��� ����/
/@/R/ d/v/4/�/�/�/�/�/ �/??�/<?*?L?r? `?�?�?�?�?�?�?�? �?O8O&O\OJO�OnO �O�O�O�O�O�O�O"_ _F_4_V_X_j_�_�_ �_�_p�_ o�_�_Bo 0ofoTo�oxo�o�o�o �o�o�o,<b P����v�� ��(��8�^�L��� p�����ʏ��ڏ܏� $��H�6�l�Z���~� ��Ɵ���؟���2�  �B�h�o������N� ԯ¯����.��R� @�v�������j�п�� ����*�<�N��^� `�rϨϖ��Ϻ����� ��$�J�8�n�\ߒ� �߶ߤ���������� 4�"�X�F�|�j��� �����������$�6� ��V�x�f��������� ������,>��N�Pb����  9� � �����$TBJOP�_GRP 2W���� ?�/��C�	�E�� � �X��X��y��^, �,{�� @� �?���D|� ��CQffC�sq3���������L���<R���D�3��[�ͨA� p��'/2'D��C&C����d/�;͟�D'�BȦ H/�/B/T/v/��/�/?333�f/ffBܦ \�/O?O  C� e5�-��/ ,2-1��?�6;����CA�f?�&ff?��CR� �R?�?b?t?��<O'J;�>y�250!+B B$cO�?��?�MAMA1E�O�F=G2j�21E�1>� �rO�O�X_B74_ _,_Z_�_f_ _�_�_ �_�_�_o�_�_:oTo�>oLozo�o~D��P��a�	V3.0�01m9a�D	*�`����%z� F&h F�C� FcP F߂� F�&p�F� F�v F��� F�� G�� G< G$� G,� G;�� GK� G\f� Gm� G�� G� G��� q�F�@ {G�pj` G�q��P G�` H�� H�pH/�� HCP HV�w =� ��
�lUn� �� (@jvT���
�?�p��oK�y� `�\�n����G����ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤߪ y�� �߬߮ !p���(�:� ��^�p����� 	������j�)���� �u�?����������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O���߳O ��S��O__�O�OK_ ]_o_�_�_�_��_�� ��_1�Y�#og�y�ko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i��O �O���O7_տ����� Ϳ/�A�S�e�wω��_����_�_�����$T�CPPACTSW�  e����IR �e�#�B�H  �SPEE/D 2� C�e��  �WwD�����_CFG K	2�#Ѵ����!Ү��_SPD��
�>�2 ���#�:�o��p�������NUM������
��OUT ;2��
  ����F����Bӳ�n�C<���z���I��������	�8���r�D�B�q��$�3�%�ZERO���  G��F�E?STPARS�#��>�F�HR��ABL/E 1����j�����t�t�t��t��Ѯ�t�	t�
Bt�t��t�t�qt�4���RDI��<�&8J\�O����$0��S��� �
� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?�����z� u���Wi{�`����n2/� 2�P`�0 3�4����2�A@��`��IMEBF_T�T���5��&ќCVE�R2�!ѯF�ќ@R �1�8�  涤 ��H7a�6����O#ѿ�� DP� [°�,_aQ|?� ��[��\_�YQ�	; '	��0[Ĕ_�Y�%�{~P��^ż�_iK<�~P��0[�oJk.a.b[1�<oNo`o�to���y
0X!�Q��$_�h�7�`_��o��ana�oVˬo��0-J�!�d` 
f���Gr��d<R�T�� !f�d�R��fu5B�rV����lis�rV�4���500P��V�l��ul�WҌ��������ÏS�`܏�o �n���0��B�T�X�h�z���1�����ğY$؟������"�4�YjH�Z�l��������cY���ʯܯ�����(�:�L�� k�c�u�����j��D�.�!�@�� �MI__CHAN�G 
̿DBGLVL�G���F��ETHER_AD ?��i�m���0r�:eu��4:3{�5:49E r�a��jqs�cP��RP��@!��!�������SNMA�SK^���o�255.$Շ�}@$�6��H�!�OOLOFS�_DI���L�OR�QCTRL D�ɦ3�:��5�T�� ������0�B�T�f� x����������������;�*�_���PE_DETAI<���֦�PGL_CONFIG WI�gA�?/cel�l/$CID$/ogrp1c�?�c�������e���2 (]o���4��3���)���40ew��� <�����/ /2/ �V/h/z/�/�/�/?/ �/�/�/
??.?�/�/ d?v?�?�?�?�?9V�e}S?�?OO*O<ONOG  O�uOTN�R? �O�O�O�O�O_L?)_ ;_M___q_�__�_�_ �_�_�_oo�_7oIo [omoo�o o�o�o�o �o�o�o3EWi {��.���� ���A�S�e�w��� ��*���я����� +���O�a�s������� 8�͟ߟ���'��� K�]�o�������������User �View ��}}�1234567890�����0�B�0J�Ӱ��j���ΩK	��?����Ͽ���  e�w�բ�	��_�qσ� �ϧϹ��*�ԣSN� �%�7�I�[�m�����ԣ5�ϼ���������u�7�}�6��p������)���}�7 _�$�6�H�Z�l�~�����}�8�������� 2��SY �lCamera٪���������E�.@毀Zl~�����  r���//(/:/ L/^/�/�/�/��/@�/�/ ??$?K�r Bɻ/p?�?�?�?�?�? q/�? OO]?6OHOZO lO~O�O7?I7��'O�O �O __$_6_�?Z_l_ ~_�O�_�_�_�_�_�_ �OI7��_Jo\ono�o �o�oK_�o�o�o7o "4FXjos^� �o�������o 2�D�V��z������� ԏ{I7�k� �2� D�V�h�z�!����� ����
��.�@�� I7��ן������¯ԯ 母�
��.�y�R�d�@v�������S�e�98� ����#�5�G��X� }Ϗ�6�����������(�߮�	t0��Z� l�~ߐߢߴ�[����� �ߣ� �2�D�V�h�z� !�3�y {������� 	��-���Q�c�u��� ��������������t ���?Qcu�� @����,) ;M_@�S;�� ����/�)/;/ M/�q/�/�/�/�/�/ r��Kb/?)?;?M? _?q?/�?�?�??�? �?OO%O7O�/�+k �?�O�O�O�O�O�O�? __%_pOI_[_m__ �_�_JO��{:_�_o o%o7oIo�Omoo�o �_�o�o�o�o�o�]  �Y>Pb t���������   Bۛ�#B������@<��B��BJU �]>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� ��2�D�V�h�z�(x  }
�`(  �2p( 	 ������ �ο��(��8�:πLς�pϦϔ��ϐ�z �^o�!�3� �oW�i�{ߍߟ߱߸S ��������F�#�5�G� Y�k�}��ߡ����� ������1�C���g� y�������������� 	P�b�?Qc��� �����( )pM_q��� ����6/%/7/ I/[/m/���/�/�/ /�/�/?!?3?E?�/ i?{?�?�/�?�?�?�? �?OR?/OAOSO�?wO �O�O�O�O�OO*O_ _+_rOO_a_s_�_�_ �_�O�_�_�_8_o'o 9oKo]ooo�_�o�o�o �_�o�o�o#5|o �ok}��o��� ���T1�C�U�� y���������ӏ��� 	��b�?�Q�c�u���8������@ ��ȟ�ڟ쟻������)frh:\tp�gl\robot�s\m900ia�&�_350_ic.xml��P�b�t� ��������ί����� �dummy "�;�?�Q�c�u����� ����Ͽ��
��.� ;�M�_�qσϕϧϹ� ��������*�7�I� [�m�ߑߣߵ������������)�;�M� _�q��������� �����%�7�I�[�m� ��������������� !3EWi{� ������� /ASew���п���;� ��88�?��"/�/@/B/ T/v/�/�/�/�/�/�/ ?�/?B?,?N?x?b?��?�?�;�$TPG�L_OUTPUT� ��  ?O�� �3;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�3 ��@2345678901�_�_�_�_ o o(c0��_Ooaoso �o�o�oAo�o�o�o'�j}1Yk} ��9K���� �1��?�g�y����� ��G������	��-� ŏ׏c�u��������� U�˟���)�;�ӟ I�q���������Q�c� ���%�7�I��W� �������ǿ_�տ�� �!�3�E�ݿ�{ύ� �ϱ�����m����� /�A�S���a߉ߛ߭�����i�A}!�� +�=�O�a�r�@/�����* ( 	 �_�������%�� I�7�Y�[�m������� ��������E3 iW�{���� ��/�V� " 7ewS���� ��RP
//�@/R/ 0/v/�/��/�/`/�/ �/�/�/*?<?�/`?r? ?�?�?�?�?�?H?�? O�?OJO\O:O�O�O �?�O�OjO�O�O�O"_ 4_�O _j_|__�_�_ �_�_�_R_oo�_Bo To2odo�o�_o�o�o to�o�o,>�ob t�����J \�(��L�^�<��� �����ʏl�ڏ �ޏ ��6�H���l�~� ��� ����؟�T��� � �V�h�F������¯ ԯv���
��.�@��� ,�v���*��������������$TPOF?F_LIM K|оӱ�|���N_SV�  �y�%� �P_�MON C�G�*�|�2y��S�TRTCHK �CE��M�VT?COMPAT:����I�VWVAR eZ���h��ϩ ��|�m��_�DEFPROG �%��%FOL�GE011ߢ�_DISPLAY����/�INST_M�SK  �� ~k�INUSER���q�LCK�܊�QU?ICKMEN��q�oSCRE�C~��tpscqԠ��!�&�%�7�_;�S�T��E�RACE_�CFG Z�����	�
?�~��HNL 2��#���� ����� ���"�4�F�X�j���ITEM 2��� �%$1234567890����  =<��������  !�����Jӫ�k��� ��);_ �/U����	 �7�	//?/ ���A/��/�/�/ 3/�/W/i/{/�/M?�/ q?�?�/�???�?A? Oe?%O7O�?MO�?O �O�?�OO�O�O�OaO 	_�O�O�O#_�Oy_�_ �__�_9_K_]_�_�_ �_Soeo�_qo�_�_�o #o�oGo}o/�o �o|�o��o��S CUg����[� ��������-�?��� c��5�G���S�Ϗ� �w�ş)����_�� ����^���y�ݟ���� �ů7����m�-��� =�c�u�ٯ�����!� ��E���)ύ�Mϱ� ÿտY�q������A� ��e�w�@ߛ�[߿�߀���ϧ��+��߀�S����F��  u�F� ��P�G�
 ]��j��(�UD1:\������R_GRP �1 ��� 	 @P������1� �U�C�y�g��������s����������?�  )I7 m[����� ��3!WEg�	�ա�q�� m�/�'//7/]/�� �/���/���/�k �/#??G?5?k?Y?�? }?�?�?�?�?�?O�? 1OOAO���O��O e/�O�O�O	_�O-_k/ Q_�/x_�/u_�_QO�_ MO�_�_oo'oMo;o qo_o�o�o�o�o�o�o �o7uOSe#_ �_������ M_3��_Z��_~��_�� ��ՏÏ����� A�/�Q�S�e������� ���џ�Eo5�G�~�SCB 2!� �����������ϯ������X_�SCREEN 1�"��
 �}i�pnl/X�gen.htm$�w����������P�Pan�el setup�ü}	index.STMÿ��1��C�U�̷
Robo�t Info e �9�ϱ��������� �τ�1�C�U�g� yߋ�߯�&������� 	��-�߶�c�u�� ����4�b�X��� )�;�M�_������� ��������x���7 I[m�6, ���!3�W�3�UALRM_M_SG ?D��Q� RD���� ��/
//:/@/q/�d/�/�/�/mSEV7  {�&kECFG $e��  E7�A1 O  B�3Q�0��492@�.�U'3rv2?D2�J?D2��b=Bn��X���b=A��Q��R�z>k�IR��X�b?+jF0h�?�2k�?�2e�d?F0�r�!GRP 2%�e� 0����Կʸ���n==�.ܽ®AcOt���OjO�O�O�O�OdI_DEFPROw�+F� (%U�P021 20 �.(_-Q0034 � %VW_USER�OD%�/_j_ �_�_�_�_�_�_o!o�oEo�GINJR �]�ONoI_MENHIST 1&e�  ( P���)/SOFT�PART/GEN�LINK?cur�rent=menupage,1�`�,2�o�o"4~��'�o�n98,1 �mp-_9U07,13�4��Dp(H�n381mp�a9����/�:��j7�q01�2mp}�������B�-�P��eedit�bFOLGE125{���"�4�?�Տ�~�p ,47  �������h�Z�\}3��20��@�*�<�G�ݟc�4�q 1,�������Ы�6a�a6o��� �2� D�V�̓므������� ȿڿi����"�4�F� X��|ώϠϲ����� e�w���0�B�T�f� �ϊߜ߮�������s� ��,�>�P�b���� ����������ݯ� (�:�L�^�p������ �������� ��$6 HZl~��� ����2DV hz����� �
/�./@/R/d/v/ �/�/)/�/�/�/�/? ?�<?N?`?r?�?�? �?�/�?�?�?OO&O �?JO\OnO�O�O�O3O �O�O�O�O_"_4_�O X_j_|_�_�_�_A_�_ �_�_oo0o�_Tofo xo�o�o�o�oOo�o�o ,>)?�ot� �����o��� (�:�L��p������� ��ʏY�k� ��$�6� H�Z��~�������Ɵ ؟g���� �2�D�V� ���������¯ԯ� u�
��.�@�R�d�Oz��$UI_PAN�EDATA 1(�������  	�}�/frh/cgt�p/respo1�.stm?_BU�SY=TRUE �=Save&AC�TION=101&C2=8p������ )prim�<�  }?�c�u�0�ϙϫϽ� )���� �����+�=�$�a�H� �ߗ�~߻ߢ���������Mv�� �5� $-$|MĨ�vagmn��� m 234&a_ctionӰ0��}�����  ual����O� ��$�6� H�Z��~�e������� ��������2V@=z�s�#� �� ������,> P�t����� ��Y/(//L/3/ p/�/i/�/�/�/�/�/  ?�/$??H?Z?�� �?�?�?�?�?�?=?O �2ODOVOhOzO�O�O O�O�O�O�O
___ @_'_d_v_]_�_�_�_ �_�_�_g?y?*o<oNo `oro�o�_�o�o-O�o �o&8�o\C ��y����� ��4�F�-�j�Q��� oo�o֏����� 0���T��ox������� ��ҟ9�����,�� P�b�I���m�����ί �ǯ��(�:����� p���������ʿ�� a��$�6�H�Z�l�~� 忢ω��ϭ�������  ��D�V�=�z�aߞ� �ߗ���G�Y�
��.� @�R�d�߈��Ͼ� ���������<�#� `�r�Y���}������� ����&J1n����}����� )�7��& cu����$� �/��;/"/_/F/ �/�/|/�/�/�/�/�/�?�������$UI�_POSTYPE�  ���� 	 �� �?��E2QUICK�MEN  T;�c3�?<RESTO�RE 1)��=i0�?��!�?�3�?��mODO VOhOzO�O/O�O�O�O �O�O�O_._@_R_d_ Oq_�_�__�_�_�_ oo�_<oNo`oro�o �o9o�o�o�o�o�_ !3�on��� �Y����"�� F�X�j�|���9C��� ��1����0�B�T� ��x���������c�� ����,�׏9�K�]� ϟ������ί௃�� �(�:�L�^������𦿸�ʿ�7SCRE��0?�=uw1sc�0u2�U3�4�5�6��7�8�E2USE1R����ks�f�U3f�4f�5f�6f��7f�8f�E0NDO_CFG *T;�g3E0PDATE� P��K�S_24�1G�_I�NFO 1+������10%  OLGGE1���� � 5�G�*�k�}�`ߡ߄� ���ߺ������1���U�g�9��OFFS_ET .�=q� l��0s���������� �!�N�E�W���[��� ����������/y��?{
j�}��UFRAME  �e�����RTO?L_ABRT�����ENB��GR�P 1/�9�1Cz  A�:8l�@8J\n������
�0Uf1�MSK  ���	-N�%��%KH/ކ2VCCM��0l��]"MR 26T9� e���f0	�g0m2%~XC5G6 *�/�&X�f4ve4�5f0A@�up��L. �8?e�7?I?v?�!hq?�?5�A�l���?�?l�� B����1l��5�?Ob??O OcONO�OrO�O�O�O �O8O�O___M_ O q_�_e���!�/�_�/ �/�/??'?o�O\o So1_�o�o�?�?�o�? __�o"io{o=jU �y���-�� �	�B�U_f�x���� �!�_���_�_�_oo 'o��\�S�1����� �o�oڟ�o_���"�i� {�=�j�U���y����� ֯-���ɯ�	�B�U� f�x����=�����͏ ߏ���'���\� S�1��ϤϷ�ɟ��� _���"�i�{�=�j�U� ��y߲ߝ���-����߀�	�B�U�f�x�O/I�SIONTMOU4� $r%���d#�7�F��G��/ FR:�\��\DATA\��� �� M�C��LOG��  � UD1��EX���' B@ ��O� �7/m�� �q���� ��  =	 1-� n6  -��U�L�&,�����O=�����U��}�TRAIN6�Ы����"8�+ (:���S.�Sas ��������'9KX&LEX�E��9�+�1-e�R,MPHASE � k%��R]!S�HIFTMENU� 1:�+
 <0\�6//�����!/ Z/1/C/�/g/y/�/�/ �/�/?�/�/D??-?�z?Q?	LIVE�/SNAPn3vsfliv��?^3}�� SETU�0�2menu�?�?d?`)O;OB��;����	(H'O�O\���Z�� ��@�A�+B8`�`��������A�B��C��G 3��KSFME�0��l��� �MO��<��z��WAITDINEND����Q@WOK  ��X[]��w_S�_^YT�IM�����\G H_�]j_�[�_�Z�_�Z<�_\XRELE�g�U@T����AS_GACT�0
h�a�鱜�d�� =��b%�$FOLGE01s1.	r000��<b�dRDIS�0�o~APV_AXSRG`2>bJ<��O��Gp~4 _IR  � �᥀������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2��D�V�h�z�����ZA�BC31?bI�� 	,�=�2��ܬ¯������
��Y���MPCF_G 1@S}0A�������ҿ�������,�b�MP��A�bI  �@���8:��Q8|O��0��t��Ϙ�?�T��� ����D����k�-ߞ����ѿp��������� ��	�l�E��i�{�� ��R�\�n߀ߚ���� ��2���e�w���� ������.��d�= OZ�s�@��\� ����'9���� Tf�����& �/5/�\// �/B/T/f/x/�/�/F ��(?:?L?v>��u��(PBS{j�P_CY�LINDER 2�CS{ ��& ,(  *�?�=�#`�?O�?8OM �/ nO�O�N�?�O$O�O�O �O_RO3_E_W_�O{_ _�O�_�_�_�_*_oof�R�2DSw�`�P�"�hoxl�s�/�o�o��o��o�o�1�qA��o*yo�o`�o� �o}�	��?y &�uJ��Z����m� ���?��׏�_�4��F����2SPHER/E 2E�=�o_�� �_��͟����_L�'� 9�i_]���⟓�z��� ������F�X�5��� Y�@�R���֯��ſ׿�N�ZZ  �$��4