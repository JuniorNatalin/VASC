��  IL�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���S�BR_T   �| 	$SVMT�R_ID $R�OBOT9$GRP_NUM<AXISQ6K 6�NFF3 _PA�RAMF	$�  ,$MD �SPD_LIT U�&2*� �� ����$$�CLASS  ������ � ��$'  1 ���  T����M-900iA�/350���aiS30/4�000 160A���
H1 DS�P1-S1��	�P01.03,�  	�  }��Pab~`�������
=�	��Xr9  ����:��D 8H�B  ������ ���  � Š���������3?����=���5w�m�c	���k��  ��/�� g���S%/� �F�� ����&Q���� ����RB� �S K ��f ��	� :?�O���'b��'/�/�/�/�/���/�/�#?5?G?Y? k?}?�?�?:� �$4*<2@2�HZl�����������8�}��c�ʘ�@m�,߈�	`��N�u C��`��4"R��<�����7�� �-#�H��� ����� B$v�?������m>'S�����P��d�T( `#� H }�� ��v$	=~'�@��OU_g_y_�_�/�_��!/�_�_� oo$o6oHoZo I��?�?63@�BOO(K��8G�y�DOVO�@lO�~O�M8� "���8�6����|�Xk��j ���� �,$�\o����#>'	Z��	����T'_*_<_��)� ;��__��_p��������ˏݏ���no�o �&12�c4�3;4@4�o�m �l�q�ٶ��2��h��~��$0��s�� (H� ��	`��/�� �6���`�����, �pRr$�'�4$B�%>!���[���.N��w.b" 6j#���v#8�yyO�ůׯ�0��V����f(�M��_�q���������˿I�(�L�65@�5p������P8G�yR��Ɵ��ܑ{�L�� �������%�@���� U$�������L�.f�(���d����7O���"���� ��u߇ߙ߫����*� ����)�;�M�_�q�&����6�6@6(�:�L��@��hBl�~ϰ�ܑ����w�ϸρ�|����G 
��p�_� ����s� �f�9��
b��I�߲�@�R�d�-?Q c�߇�ߘ�����);�����<TqPHP�8u	u��o �����//,/ >/P/b/t/�/�/�/�/ �/�/�/?<�?8? J?\?n?�?�?�?�?�? �?�?�3n`
O�� �pO�O�O�O�O�O�O �O __$_6_H_Z_l_ ~_�_�_�_�_"?�_�_ o o2oDoVohozo�o��o�;  =��EXTENDED_ AXIS-��q���4/5�� oH h� -ND���0.33���  �PG�Tq�H�X{�~q����&��{�'�9~��5
� ���r �l3� �ܑt▂ ������ �,��cڐ� 7� (^rt Z��	�!��_�q�����3� ����ӏ���	��-�?�Q�c��(OO|� >OPObO�����*� <�N�`�r��������� ̯ޯ���&�8��_ \�n���������ȿڿ �����?����Yϴ� Ɵ�Ϡϲ��������� ��0�B�T�f�xߊ� �߮�������@��� ,�>�P�b�t���� ����*�<���`�rτ� L�^�p����������� ���� $6HZ l~������� � 2DVhz ������0�B�
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?��?�?�?�? �?�?�?OO&O8O� ���O���O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oh?0oBoTofoxo�o �o�o�o�o�o�oROdO �O�O�Ot��� ������(�:� L�^�p���������ʏ &o� ��$�6�H�Z� l�~������o0"̟ FXj2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v���� ����п�����*� <�N�`ϼ������� �������&�8�J� \�n߀ߒߤ߶����� �����"�4X�j� |������������ ��zό�6������� ������������ ,>Pbt��� ����N�(: L^p������&�  =�E�XTENDED �AXISh����aiS4/50�00 40Ak��H  DSP -�~�P00.39��� 	�  �o�Pm� H��X�q����_�  {n�C �9~�5
�? �p� �l� l����tn� b��/�/�/�/
??.?�e�c	`�� 7 (�"t �Z� :�?�j��!>?�?�?�?�?n��?�?OO'O9O`KO]OoO�O�O�X� J��On�����_$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo ho�o�o�o�o�o�o �o
.@,��O�O ��O�O����� �*�<�N�`�r����� ����̏ޏ����po 8�J�\�n��������� ȟڟ���Zl�� ��|�������į֯ �����0�B�T�f� x���������ҿ.��� ��,�>�P�b�tφ� �Ϫ���*i!/%/ 7/I/[/m//�/�/�� �߸������� ��E? W?i?{?l�~����? ��������� �2�D� V�h��O=�/���S�e� ����	-?Qc u������� );߿Mq� ������// %/���=/�������/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?UO/OAOSO eOwO�O�O�O�O�O-/ _/Q/�Ou/�/�/a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�oO�o�o�o# 5GYk}��O_ _�3_E_��1�C� U�g�y���������ӏ ���	��-�?�Q�c� �ou�������ϟ�� ��)�;�M���e� ���˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�}� E�W�i�{ύϟϱ��� ������U���y�#ߝ� �����ߛ߭߿����� ����+�=�O�a�s� ���������;�� �'�9�K�]�o����� �����E�7� [�m� 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�����/+�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO�mOO�O�O �O�O�O�O�O_!_}/ �/�/K_�/�/�/�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �ocO+=Oas ������;_m_ __(��_�_]�o����� ����ɏۏ����#� 5�G�Y�k�}������� ş�����1�C� U�g�y��������� /�A�S��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�q�͟ �ϧϹ��������� %�7�Iߥ�ׯɯs�� ����������!�3� E�W�i�{������ ��������/���S� e�w������������� ��cߕ߇�P�߽� ������� '9K]o�� ����7��/#/ 5/G/Y/k/}/�/�/�/ �/!3�/Wi{C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O��O�O�O�O __)_;_M___q_�/ �/�/�_?'?9?oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EW�O{���� �����/��_�_ �_x��_�_����я� ����+�=�O�a�s� ��������͟ߟ�� _�9�K�]�o����� ����ɯۯ�I�[�� �����k�}������� ſ׿�����1�C� U�g�yϋϝϯ���� ����	��-�?�Q�c� u߇ߙ���'����=� O�a�)�;�M�_�q�� ������������ %�7�I�[�m���ϣ� ����������!3 EW�����ߠ��� ���/AS ew������ �//+/��=/a/s/ �/�/�/�/�/�/�/? ?q�-?����? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�OE/__1_C_ U_g_y_�_�_�_�_? O?A?�_e?w?�?Qoco uo�o�o�o�o�o�o�o );M_q� ��_����� %�7�I�[�m���_o �_ȏ#o5o���!�3� E�W�i�{�������ß ՟�����/�A�S� �e���������ѯ� ����+�=�����U� Ϗ�󏻿Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������m� 5�G�Y�k�}ߏߡ߳� ������E�w�i� ����y�������� ����	��-�?�Q�c� u�����������+��� );M_q� ���5�'��K�]� %7I[m�� �����/!/3/ E/W/i/{/���/�/�/ �/�/�/??/?A?S? e?��}?�	�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_�/]_o_�_�_ �_�_�_�_�_�_om? �?�?;o�?�?�?�o�o �o�o�o�o1C Ugy����� ��S_�-�?�Q�c� u���������Ϗ+o]o Oo�so�oM�_�q��� ������˟ݟ��� %�7�I�[�m������ ���ٯ����!�3� E�W�i�{�������� �1�C���/�A�S� e�wωϛϭϿ����� ����+�=�O�a߽� �ߗߩ߻�������� �'�9ǿ��c�ݿ �����������#� 5�G�Y�k�}������� ��������{�C Ugy����� ��S��w�@��� u������� //)/;/M/_/q/�/ �/�/�/�/'�/?? %?7?I?[?m??�?�? �?#�?GYk3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�/�_�_�_�_ �_oo+o=oOoao�? �?�?�oOO)O�o '9K]o�� �������#� 5�G��_k�}������� ŏ׏�����{o�o �oh��o�o������ӟ ���	��-�?�Q�c� u���������ϯ�� O��)�;�M�_�q��� ������˿ݿ9�K��� o�����[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱�� ��������/�A�S� e�w����	ϳ�-� ?�Q��+�=�O�a�s� �������������� '9K]o�ߓ ������# 5G���������� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??w-?Q?c? u?�?�?�?�?�?�?�? OasO����O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_5?�_o!o3o EoWoio{o�o�o�oO ?O1O�oUOgOyOAS ew������ ���+�=�O�a�s� �����_��͏ߏ�� �'�9�K�]�o��o�o �o��%����#� 5�G�Y�k�}������� ůׯ�����1�C� ��U�y���������ӿ ���	��-ω���E� ��џ㟫Ͻ������� ��)�;�M�_�q߃� �ߧ߹��������]� %�7�I�[�m���� ������5�g�Y��}� �ϡ�i�{��������� ������/AS ew������ �+=Oas ����%���;�M� /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?�}?�?�? �?�?�?�?OO1OCO UO��mO��/�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo)o�?Mo_oqo�o �o�o�o�o�o�o]O �O�O+�O�O�O�� ������!�3� E�W�i�{�������Ï Տ�Co��/�A�S� e�w���������M ?�cu=�O�a�s� ��������ͯ߯�� �'�9�K�]�o����� �ɿۿ����#� 5�G�Y�k�}�ٟ럕� �!�3�����1�C� U�g�yߋߝ߯����� ����	��-�?�Qﭿ u����������� ��)��Ϸϩ�S��� ���Ϲ������� %7I[m�� �����k�3 EWi{���� ��C�u�g�0/���� e/w/�/�/�/�/�/�/ �/??+?=?O?a?s? �?�?�?�?�?�?O O'O9OKO]OoO�O�O �O//�O7/I/[/#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCo Uogoyo�?�o�o�o�o �o�o	-?Q�O �O�O{�O__�� ��)�;�M�_�q��� ������ˏݏ��� %�7��o[�m������ ��ǟٟ����k� �X���������ï կ�����/�A�S� e�w���������ѿ� ?����+�=�O�a�s� �ϗϩϻ���)�;��� _�q���K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}����� ����������1�C� U�g�y�����ϣ�� /�A�	-?Qc u������� );M_�� ������// %/7/�������/���� �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?�?�?OgOAOSO eOwO�O�O�O�O�O�O �OQ/c/_�/�/�/s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o%O�o�o# 5GYk}���O /_!_�E_W_i_1�C� U�g�y���������ӏ ���	��-�?�Q�c� u����o����ϟ�� ��)�;�M�_��� �����ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� ��E�i�{ύϟϱ��� ��������y���5� ����ӯ�߭߿����� ����+�=�O�a�s� �����������M� �'�9�K�]�o����� ������%�W�I���m� ߑ�Yk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/���/+= ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[O�mO�O�O �O�O�O�O�O_!_3_�E_�$�$SBR2� 1�%qP T0 � �/�) �_�_�_�_�_�_ oo,o>oPoboto�o �o{_�_�o�o�o (:L^p��� ��o�o�o ��$�6� H�Z�l�~�������Ə ؏����2�D�V� h�z�������ԟ� ��
����@�#�d�v� ��������Я���� �*�<�N�1�r�U��� ����̿޿���&� 8�J�\�nπ�c�L_�� ����������,�>� P�b�t߆ߘߪ߸ٚ� �������"�4�F�X� j�|��������� ����#�5� G�Y�k�}��������� ��������0BT fx������ �,>��bt �������/ /(/:/L/^/p/T�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�/ �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �?�O
__._@_R_d_ v_�_�_�_�_�_�_�_ o�O*o<oNo`oro�o �o�o�o�o�o�o &
oo\n��� ������"�4� F�X�<h�������ď ֏�����0�B�T� f�x���n�����ҟ� ����,�>�P�b�t� ������������� �)�;�M�_�q����� ����˿ݿ�"�$� 6�H�Z�l�~ϐϢϴ� ��������� ߤ�D� V�h�zߌߞ߰����� ����
��.�@�R�6� v����������� ��*�<�N�`�r��� د���������� '9K]o��� �j����"4 FXj|���� ����//0/B/T/ f/x/�/�/�/�/�/�/ �/?�?>?P?b?t? �?�?�?�?�?�?�?O O(O:O?^OpO�O�O �O�O�O�O�O __$_ 6_H_Z_l_PO�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�_�o�o �o�o
.@Rd v������o� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� �X�j�|�������į ֯�����0�B�T� f�J���������ҿ� ����,�>�P�b�t� ��j�|���������� �(�:�L�^�p߂ߔ� �߸ߜ����� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
 �@Rd v������� *<N2r� ������// &/8/J/\/n/�/d�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�/ �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �?__,_>_P_b_t_ �_�_�_�_�_�_�_o o�O:oLo^opo�o�o �o�o�o�o�o $ 6o,ol~��� ����� �2�D� V�h�Lx�����ԏ ���
��.�@�R�d� v�����~���П��� ��*�<�N�`�r��� ������̯����� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0��T� f�xߊߜ߮������� ����,�>�P�b�F� ������������ �(�:�L�^�p����� x�������� $ 6HZl~��� ����� 2D Vhz����� ���/./@/R/d/ v/�/�/�/�/�/�/�/ ??�(?N?`?r?�? �?�?�?�?�?�?OO &O8OJO.?nO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_`O�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�_�o�o �o,>Pbt �������o� �(�:�L�^�p����� ����ʏ܏� ��� 6�H�Z�l�~������� Ɵ؟���� �2�D� (�h�z�������¯ԯ ���
��.�@�R�d� v�Z�������п��� ��*�<�N�`�rτ� ��z����������� &�8�J�\�n߀ߒߤ� ���߬������"�4� F�X�j�|������ ���������0�B�T� f�x������������� ��,�Pbt ������� (:L^B�� ����� //$/ 6/H/Z/l/~/�/t�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�/ �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O �?_*_<_N_`_r_�_ �_�_�_�_�_�_oo &o
_Jo\ono�o�o�o �o�o�o�o�o"4 F*o<o|���� �����0�B�T� f�x�\������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ�� ��$� 6�H�Z�l�~������� ƿؿ�����2�D� V�h�zόϞϰ����� ����
��.�@�$�d� v߈ߚ߬߾������� ��*�<�N�`�r�V� ������������ &�8�J�\�n������� ����������"4 FXj|���� ����0BT fx������ ���,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?/8?^?p?�?�? �?�?�?�?�? OO$O 6OHOZO>?~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_pO�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�_�o�o *<N`r� �������o� &�8�J�\�n������� ��ȏڏ����"�4�