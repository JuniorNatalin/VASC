��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �
  ����
��WVAMP_T �  $X�1  $X2�AY@.�/FC~5  $2�ENBA $DTo  / _R2� d ENAB�LEDnSCHDo_NUMA  x�CFG5� $GROUP�}$z ACCEL@��G$MAX_OFREQ�2 L��DWEL�DEB�UG�PREWS�OUT�PU�LSEASHI�Ft 7TYP4�$USE_AEF|} 4$GDO��  f0 �r?�NpWEA�VE_TSK ��V�_GP�S�UPPORT_C�FnCNVT_DONE p }k�}GRP 2�r�� _� �$>� TIME1�o:$2'EXT� (�1#&(MODE_S�W�CO3 SWI�T � �/ PHA|X6  4 � �ECC$�TE�RMNnPEA�Kno!AL O \ � �!I�k$�!N_VSTAR�#!r"���"�%�CYCmL42 �/ �� Tv"b $CUR_REL_� �! �/ WPR�5 � 
$C�EN� _RI3R�ADIU�X�Iz ] ZIM�UTi!$ELE?VATIONg5� �N�CONTIN�UOe2q �MEX�AC=PE��81�6  H~ ��UENCYA�I�TUD4�2RIG�HC�2LEBL_�ANG1 �O�TF_� 	��  $3A�bE�T��n3C!�$ORGjHFB)KjH��P��C�.�DLDW�HR�E�_�3�B�C��D�B�Cp�@�D�A�CCHG�G�	Q�F	Q�F	Q�FINC�G=Q�F=Q�F=Q�F؃AVCPYC� _T��\#�Y~P#�@SY��H)@�UPD�"0n�$$CL�ASS  �C���Q��8 �P�� �VA2�Uw� � ?��@�  aa�U�T o-o?oQoco�P�TNw 2 �[ f���ue@O߀i�oc�Q� � �Ua	`��`�d �`� �����=�������b  ����.pqUcw-� ut(q��uvp�P��x u��d�aPq�&��8���
�s,��}a� u s�s�a�s��������֏b�Q�  2��[
TacSI��}�v��F�j ,�?1�'�� P�0��P�P�a��0� l�jk��ҟ������,�>�llFI�GURE 8�� 3�:�a0�*�X�e�ۯ ү�������L�R��d�v������T'CIR1q�dֿ A���B�,�>���0�����:�`�B��ϲ�p������nj�� pq�(qG�V�E�@ �����`+ݳ��ߗ� �߻���������'�<9�S�L��%��B�5)��T�` ���p���䏟��w� �#�5�G�Y�k�}����mkTrianglej���>�,� ��L���D�Qcu�������� �������X�+X 2D�����/ /'/9/�},> l/�/���/?!?�3?E?W?i?{?�?�� C��?nhE��?�?O O,O>OPObOtO�O�O �O�O�O�O�K�?�O�? �?H_Z_l_~_�_�_�_ �_�_�_�_o o2o|m�SCHEXTEN�B  ��c�STATE 2�k @o�o�o�o�o~NgWPR ����}��_OTF' 	�oa�@� qq�]qQcuv�quA��os�u@�  <#��
�?��^�1u_�GP 2;| � Io(�:������ ��e+