��   v��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<�$1_8k ���FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\9 ^75z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D`�VCAX_�w A.  @ 5vFX0OR�@E ?NUM_SE238�_TO0Q�#RE_:� 2cT �+V>1 , $� �ME�vUPgDAT�wAXy_2 	�+VS5Q' 8<P��PnP;0k L\�R�PA�kQ�Q��+VM5Q  �$ISRTd 5+VG5Q { v��R2 
v�S2�T kR9�P 	��$U1SS  O����a����w�$' 1 �e� } �� 	 ����o�o�o�e�����
������L) ����2����b�`���31V��3��g��or�
p�Jp�t�~�o�t��o�c�K}�����d ��7{`�P�&�.�`����|��+�=�d�a�A����� � :Z�  �����w�B ��  䲁�`f�p���������K��_������.��J~��l���j���.���_N �/�2���d�1�xC�U���=L��`�f��?�����@��� ͟ߟ���'�9�K�`]�o������� �eྯ̧��쯄d  2  ��/�A�S�e�w�����������<���� ��1�C�U�g�yϋ� �ϯ����`�a�o��� ���*�<�#�`�K߄� oߨߓ�c��ߡ���� &�[�5�G�n�k�}�� �����������"�� �P�b�t��������� ������(:�� ^p������E ϯ��6HZl ~�����˿� / /2/D/V/h/z/�/ �/�/�/�/���/��/ .??R?9?v?a?�?�? �?�?���?�?OO<O 'O�?]OoO�O�O�O�O 3O�O�O_�O_J_=� k_}_�_�_�_�_�_�_ �_oo1oCoUo|o �o�o�o�o�o�goio �o-#Tfx�� �������,� >�P�b�t��������� Ώ����/�(��L� 7�p�W������ʟ�� ��?�՟6�!�Z�l� �O{�������ïկQ� ���2�D�/�h�[_�� ������ѿ����� +�=�O�a�s�5�Ϭ� ��������G���'� K�Ar߄ߖߨߺ��� �������m�J�\� n�����������������$FMS_GRP 1^�� �>�J
�H �C?H�-�I����J��I��X�J�Mb.�O��OL� K�1�UJ(H�J��qJ�B�  ����BV'B���9B����²Z�B���8J����u��U�|PD�O����K��nJ��ߘK
X���=��?���J
�WH I�H�1�4I���J�	�I�Y�+�VBP����V����������3� �� ���  	Q�+j;nQSJ_�QSK� ���OC�OC�WW-OPyC�O�m P/�&�k.kAP��w7w<Q�P�;GX�%X�+8�4����&�8���i�������p���S������.�������h	��9�����������y.Y��p����P���g���i��H���G^�� /����_7%�^�%�����ݟ��G����������2���+�� �?��w���_{�N���j~�w9��vk����%��7 ��� ���������k� ��O �� "��g "�� "k�X "Nv ���5 ������#��n����?��(Z��?��� � � ���0"�o4��yV��g��r;]4��]5�e�C�e��e���e��{��h�a�%���,���z�Zz��� �sHq�g�7��>�����f&��<�V��� h�����l�r'0���l�I/0����$E�s*T�������*������NK0*���M��������"6�Y�;��Y����'���=�������0�`���c��d��0��uA��W�Y�:���/��Ւ�	�t�0��2
����Z	Ec"}��;
P�4�=�?�?d�4C4�}!_������
��D�4�0�  ?���uN
��P�	��"_�l_�s4��74�,(�V��?,���VJ�V	�
�,��[D�_ФJ4��@%��$
�}'� �  �i	+�_�����Y[DU�_��@�� �
��	��{H$@�����I�	����_�[D�_Л$@��$@&�_���	����P��nURQ�ī��4R4�K@��$@(��E��+�����@�V�X��4eoo'o9o?b�3Yo FVvo�o�4�U�d>�E4�1�dS�l�a�1z�h�i�a�7>k��>k�˰?L9?H��:?o!�?o�?l��?m��?mE3?m��W>I8&>^��O?j��?j��u?j�v?j��p;s��?j��~>l�<7=��uv=�/�>���?)?�*F?�?)�Ai?)F�?)�Ot?)X�<��񼼝?��m?��?
�S+?	�ʏp���pj?�=��iZ7���J���'��Ĵg��̧��������,��cֿ��k���x����1���@�������]����x����a���D��t_����2��uC7<����<�q�?���@ �?���e?��F?��B_?�A�?��E ?�;!����ּ;�6?��n\?�I�?��\?��6�3?���<�)a7������ϻ������-���8._������tg�v�ӓ���ӖV�������ne������#���㘯��6K��J��u���	'��~���b�� >�����W�F�_��?�k�?�b�?���?����?���?���>�j>��?� �?��	�?�}�?����߄�?�|>��	,($UP00�a �'���4���X�?�USER_ADVi�k�Q�����ޟ�ŝMAKRO080���>�%�b�I� [���ϟ������򯁯 ����L�3�p�W�y� {���ʿ���ͯ߯$� �H��l�W�iϢύ� �ϱ���������D� /�h�Sߌ�s߰ߛ߭� ����
��9�kY� k�}���߳���T��� �����1�C�U�g�&� ��������������	 ��-?Qc"�� ��|���) ;M_���� x��/�%/7/I/ [///�/�/�/t/�/ �/�/�/!?3?E?W?? {?�?�?n�Rp?�?�? �?d?O/OAOSOOwO �O�O�OlO�O�O�O�O _+_=_O__s_�_�_��_h_�_�_�_�[��1�234567890o'eu�oIo9omo ]oyo�o�o�o�o�o�o �o!-5G{k �������� ��S�C�_�g�y��� ������ӏ����� 7�a���ﲟ�� �ӟ���0��T�?� x�c�u�����ү���� ��,�#�P��_t��� ����	����o��� (��L�^�pς�AϦ� �����ϛ� ��$��� H�Z�l�~�=ߢߴ��� �ߗ���� ���D�V� h�z�9�������� ��
����@�R�d�v� 5������������� ��<N`r1� ���?�� 8J\n-��� ����/�4/F/ X/j/)/�/�/�/�/�/ �/�/?oc�9?Q�]? M?i?q?�?�?�?�?�? �?OOO%O7OkO[O wOO�O�O�O�O�O�O �O_C_3_O_W_i_�_ �_�_�_�_�_�_oo 'oQoAouou�?�o�o �o�o�o�o D/ Aze����� ����@�7�d�v� �/������Џ/�􏃏 �*�<�N��r����� U���̟ޟ🯟�&� 8�J�	�n�����Q��� ȯگ쯫��"�4�F� �j�|���M���Ŀֿ 迧���0�B��f� xϊ�IϚ������ϣ� ��,�>���b�t߆� Eߖ߼�������� (�:��^�p��A�� ������� ��$�6� ��Z�l�~�=������� ������ 2)?M eoYas���� ��'[K go������ ��3/#/?/G/Y/�/ }/�/�/�/�/�/�/�/ ?A?1?e?U?q?y?�1��$PLCL_G?RP 1���1�� �D�0�?�  ��:`?t�� �9�O�:O%O^OIO �OmOO�O�O�O�O _ �O�>2_�OY_�O}_h_ �_�_�_�_�_�_�_o 
oCo*o$_vo8o�o4o �o�o�o�o	? *cN�nho�| �x��)��M�_��J���n�����ˏ=��$VCAX_RE�F�0 2�5� t �
 ���ER�ENCE 1�� ׏7�I�[�m�������2�ԟ���
��.�@����3ß|��������į֯�S��4 k�$�6�H�Z�l�~������5�̿޿�� �&�8ϣ���4��zπ�Ϟϰ������ϱ�7 c��.�@�R�d�v߈����8��������� ��0���9��l�~��������C��FACTORY DATA\��'�9�@K�]�o������9�������������	� ��GYk
�2_���������2_�P bt����'j� ?�
//./@/R/d/ '���/�/�/�/�/ �/?'���/H?Z?l? ~?�?�?�?'b�7?�? OO&O8OJO\O'
� �?�O�O�O�O�O�O_ '�ՇO@_R_d_v_�_ �_�_'Z�/_�_�_o o0oBoTo���_�o�o �o�o�o�o�o�� /ASew%�����3��%�7� I�[�m���_�t7�� Ώ�����(����� �d�v���������П ;����/��0�B�T� f�x�㟥�/?��Ưد ���� ������?\� n���������ȿ3��� O��(�:�L�^�p� ۿ��'_�Ͼ������� �߃ϥ��_T�f�x� �ߜ߮���_oqo��� �,�>�P�b�t�� ����������(�:�L����4����� ����������*�p��� 0BTfx�� S���� 2 D������� ���W��(/:/ L/^/p/�/�/�K� �/�/�/??*?<?�/ �x?�?�?�?�?�? �?O?�� O2ODOVO hOzO�O�?C��O�O �O�O_"_4_����j_ |_�_�_�_�_�_�_�� 	�o!o3oEoWoio� �o�o�o�d