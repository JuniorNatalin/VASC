A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DRYRUN_T   � $DRYRUN_ENB  $NUM_PORT  $NUM_SUB  $STATE  $TCOL_SYSPT  $PMC_SYSPT  $GRP_MASK  $STEP_MOTION  $LOG_INFO  $TCOL_SAVE  $FLTR_EMPTY  $PROD_START  $ESTOP_DSBL  $POW_RECOV  $OPR_DSBL  $SAW_PROG %$INIT_PROG %$RESUME_TYPE  ��DRYRUN_PORT_  4 $TYPE  $FST_IDX  $LST_IDX  $STATIC_PORT  ���MIX_BG_T  4 $PROG_NAME %$MODE  $STATUS  $MODIFY_TIME   �MIX_MKR_T   $LINE   $LINE_SIZE  ��MIX_LOGIC_T , $USE_FLG  $USE_MKR  $USE_TCOL  $USE_TCOLSIM  $NUM_FLG  $NUM_MKR  $NUM_BG  $NUM_SCAN  $MAXNUM_SCAN  $MINNUM_SCAN  $ITEM_COUNT  $PROC_TIME  $MAX_TMR_VAL  $TCOL_LINE $TCOL_ENB  $TCOL_SIM  $TCOL_STAT  $SAVE_IDX  $SAVE_LINE $TCOL_WARN  $BG_HITEM  $INST_CHK  �$$CLASS  ������   5    5�$DRYRUN  ������5�      c                        ����                   %VAGSAW                                %VAGTPINI                                 �$DRYRUN_PORT 2������5� c    "      $             d                   )     �                                             	  	                    �  �         �  �         �  �         �  �         �  �                    !  8         c  c         h  i         l  l         y  �         �  �         �  �         �  �                      	                      2         9  ;         A  P         a  x         �  �         �  �         �  �         �  �         �  �         �  �         �  �         �  �           !         )  +         C  C         H  I         L  L         Q  q         y  {         �  �         �  �         �  �         �  �         �  �         �  �         �  �         	  	         !  3         7  7         I  I         a  s         w  w         �  �         �  �         �  �                                 1  A         V  a         v  �       )   D   G       )   M   P       )   y   z       )             )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )           )  !  !       )  2  2       )  J  J       )  A  A       )  P  P       )  `  c       )  e  e       )  u  x       )  z  z       )  �  �       )  
  9       )  �  �       )  �  �                                                                                                    �$DRYRUN_SUB ?������5�  FOLGE         UP            MAKRO      ) SUCHL         BIN1         x�$MIX_BG 2������5�  4%MAKROSP1                                    JQ�%MAKROSP2                                    JQ�%MAKROSP3                                    ����%MAKROSP4                                    ����%MAKROSP5                                    ����%MAKROSP6                                    ����%MAKROSP7                                    ����%MAKROSP8                                    JQ��$MIX_LOGIC ������5�                  �              X  ����  s2tt* q*  q* !q
squ
tt* !qs)Sr)�tt
tt                                                                                                                                                                                                                       ����  s2tt* q*  q* !q
squ
tt* !qs)Sr)�ttqu
Kq
Lttttt�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������             �$MIX_MKR 2������5 �  * dss
]q
_q
_tr
 t                                                                                                                                                                                                                                         * dsu
]qu
_qu
`t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ds
 +q
 -q
 /q
 1t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    * ds
 q
 q
Rt                                                                                                                                                                                                                                                * ds
Cqu
Dq
Equ
Fq
Gqu
Hq
Iqu
Jq
Kqu
Ltt                                                                                                                                                                                                     =  *  dsu
Cq
Dqu
Eq
Fqu
Gq
Hqu
Iq
Jqu
Kq
Ltt                                                                                                                                                                                                     =  * !dsu
Mq
Nqu
Oq
Pt                                                                                                                                                                                                                                         * "ds
Mqu
Nq
Oqu
Pt                                                                                                                                                                                                                                         * #ds2 tOqu
Pq
Qqu
Rt                                                                                                                                                                                                                                       	  * $ds2 tOq
Pqu
Qq
Rt                                                                                                                                                                                                                                       	  * %ds2 tSqu
Tq
Uqu
Vt                                                                                                                                                                                                                                       	  * &ds2 tSq
Tqu
Uq
Vt                                                                                                                                                                                                                                       	  * 'ds2 t                                                                                                                                                                                                                                                          	  * (ds2 t                                                                                                                                                                                                                                                          	  * )ds2 t                                                                                                                                                                                                                                                          	  * *ds2 t                                                                                                                                                                                                                                                          	  * +ds2 t                                                                                                                                                                                                                                                          	  * ,ds2 t                                                                                                                                                                                                                                                          	  * -ds2 t                                                                                                                                                                                                                                                          	  * .ds2 t                                                                                                                                                                                                                                                          	  * /ds2 t                                                                                                                                                                                                                                                          	  * 0ds2 t                                                                                                                                                                                                                                                          	  * 1ds2 t                                                                                                                                                                                                                                                          	  * 2ds2 t                                                                                                                                                                                                                                                          	  * 3ds2 t                                                                                                                                                                                                                                                          	  * 4ds2 t                                                                                                                                                                                                                                                          	  * 5ds2 t                                                                                                                                                                                                                                                          	  * 6ds2 t                                                                                                                                                                                                                                                          	  * 7ds2 t                                                                                                                                                                                                                                                          	  * 8ds2 t                                                                                                                                                                                                                                                          	  * 9ds2 t                                                                                                                                                                                                                                                          	  * :ds2 t                                                                                                                                                                                                                                                          	  * ;ds2 t                                                                                                                                                                                                                                                          	  * <ds2 t                                                                                                                                                                                                                                                          	  * =ds2 t                                                                                                                                                                                                                                                          	  * >ds2 t                                                                                                                                                                                                                                                          	  * ?ds2 t                                                                                                                                                                                                                                                          	  * @ds2 t                                                                                                                                                                                                                                                          	  * Ads2 t                                                                                                                                                                                                                                                          	  * Bds2 t                                                                                                                                                                                                                                                          	  * Cds2 t                                                                                                                                                                                                                                                          	  * Dds2 t                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                _ds
�qu
�q
�q
�qssu
�q
�tr�tqu
qu
q�t                                                                                                                                                                                                        `ds
Jqu
Lqu
Kq
Mqu�qs)Arskq) �trsq) �ttt                                                                                                                                                                                                       adss
�q�r)8tq
BqBqu) Hqu) Iqs) Zr) \tt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     