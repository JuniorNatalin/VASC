��   �A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG��DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST���DwNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !���* D� $PRIMA�R_IG !$ALTERN1�<WAIT_TI|A ���FT�� @� LOG�_8	�CMO>�$DNLD_FI�:�SUBDIR�CAP� ����8 . 4� H��ADDRTY�P�H NGTH���4�z +LS��&$ROB{OT2PEER2ބ MASK4MR�U~OMGDEV�� RCM�  $Z ��QSIZ�X�� �TATUSWMA�ILSERV �$PLAN� <�$LIN<$C�LU���<$TO��P$CC�&FR\�&�JEC�!�%�ENB � ALkARl!B�TP��3�V8 S��$�VAR9M ONx
6��
6APPL
6�PA� 5B 	7PO�R��#_�!�"AL�ERT�&�2URL� }�3ATT�AC��0ERR_oTHRO�3US�9z!�800CH- Y�4�MAX?��RD�M*T $DI�S� ��SM�B�	"�BCA��$WI2A{IN4EXPS�!n�PAR��0B{CL�
 <(�C�0�SPTMOU�4� WR�_HuF� �0@o !l5��!�"%�7X�ECC�%� V�R�0UP� _DL�V�vE��SNo3 �O�BX�_S@~#Z_IND9E
B�QOFF� ~kUR�YD��KT��   t 9�!&PMON��S�D��RHOU�#E�ND�X�Q�V�Q�VL�OCA� Y$Nޅ0H_HE��OTCPI"/ 3 $ARPz&�1�F�W_\ �I!F,�P;FA~Lk01#�HO_� INF�O7cEL	% P� K  !k0WO��@ $ACC�E� LV�K�2�H#ICE��` ��$�c# ����q��
��
�$�'0 u
�*��F����ItDuw�$� 2,{T ��r|}]p�� ,}��!q����r%r,z���0�At�Dq�s`_  ,{�Krr������� ��̏ޏ����&�8���t� _FLTR � v4s ��
�������{nx,}�2�{ZbSHw@D �1,y  P��Atџ���2� ��V��z�=���a��� ԯ�������߯@�� d�'�9���]������ ���ɿۿ<���`�#� ��GϨ�kϡ������ ��&���J��V�1�� ��g��ߋ��߯���� 4���	�j�-��Q�� u��������0��� T��x�;�q�������p�����wz _LI� �1]�x!1."10����01A��255.y8���Iu/26H�  \n���3�H@%���
�4&�H�L^p��5 �H �����6/H� </N/`/r/�L�RCj`�pp�!Pp%�ː�v� Q� ���.<(?]?o? B?�?�?�?�?�?�?��P�?O/OAO OeOwO��O�OZO�O�O�O�. �O��Lu-_\_�Or_��_�_�_��}iR�Connect:� irc�T//alerts�_�_o o%o�Ul_Qocouo�o�o�o����  j�"<��d� DM%s��~�$SMB 	���@o�/C��v�`_CLNT �2
�� 4#T -�\����� ��3��$�i�H������~�ÏՏ����NM���n%�L�T��:�{��j�����Hǟ\�aN�1�m�%172.2�0� 4�3ӟ(v�������8����#�USTOM ��m3���0 ����$TCPIP��b�mX5 TKEL�e1�2��H!TP!�#{�rj3_tpd�ן # ��!K�CL�諻���)u!CRTB�0����2�!CON�S�����smo	n���