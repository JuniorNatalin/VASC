A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �SBR_T   | 	$SVMTR_ID  $ROBOT_ID $GRP_NUM  $AXIS_NUM  $MTR_ID $MTR_INF_ID $SV_PARAM_ID 	$PARAM  ,$MOT_SPD_LIM   ��SBR2_T   $PARAM   �`���$$CLASS  ������       �$SBR 1 ������ T�    R-2000iB/185L               aiSR30/3000 80A       
H1 DSP1-S1    	P01.03    ,  	�     PAR      ����   �    
=  
#�r9  ~��%�        8 l�  ���x� %        �       ��      ��   ��  2'-b��>��q�G�R����          &��� % ���� �      �                       ����        	��w��N��          �c9	`B 0     � �� :?p�   @  'bx�                                                                                                                                  3                                                            Z                 2�'{��>O�r�+� 3 ���=�����1�%m�                                          �    R-2000iB/185L               aiSR30/3000 80A       
H2 DSP1-S2    	P01.03    ,  	�     PAR�      ����   ��    
=  
8��r9  ~��%�        8 l� ,p�@� n        ��       o�o�      ��   #q 3 ���=����k)2!�h	��          &��u  ���� u      �t                       ���.        ��-k����         �c9	`B 0     � �� :?p�   @    x�                                                                                                                                  3                                                            Z                 3�2��<����n	��0�4h���<z�1�`��D	�                                          �    R-2000iB/185L               aiSR30/3000 80A       
H3 DSP1-S3    	P01.03    ,  	�     PAR�       ����   �@    
=  
3�Ir9  ~��%�        8 l� @��x� n        ��       keke      ��         2�#���>�v�l��^7
�          &�      ���� U      �V                       ���_        	b����	��M         =c9	`B 0     � �� :?p�   @    x�                                                                                                                                  3                                                            Z                                                                                                   �    R-2000iB/185L               aiS12/4000 40A        
H4 DSP1-S4    	P01.03    ,  	�     PC        �q��   2��    
=  
8��r9  ~�$0        � (H�  ������F        � �                  �                                                     0 ���� Y      ��                       ���$         ��9	b��/���         ��       �� :?�          y                                                                                                                                  f                                                                                                                                                                      R-2000iB/185L               aiS12/4000 40A        
H5 DSP1-S5    	P01.03    ,  	�     PC        �q��   2��    
=  
8��r9  ~�$0        � (H�  ���@��
         � �                  �                                                     + ���� Z      ��                       �)�I         0����Q���         ��       �� :?�          y                                                                                                                                  f                                                                                                                                                                      R-2000iB/185L               aiS12/4000 40A        
H6 DSP1-S6    	P01.03    ,  	�     PC        �q��   2�     
=  
8�r9  ~�$0        � (H�  �������       �                  �                                                     F 
���� \      ��                       �           ��4��vu�         ��       �� :?�          y                                                                                                                                  f                                                                                                                                                                  �  @�EXTENDED AXIS               aiS22/4000 160A       H  DSP -      	P00.39    ,  	�       P         E����   �z��  {      r    ��9 :    � 8H	�         ���                                                                                                                               }            %p�                    B	�  P     c Z� :?��          �                                                                                                9                                                                                                                                                                                                      �����                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  =�EXTENDED AXIS               aiS4/5000 40A         H  DSP -      	P00.39    ,  	�       P         H�X�   ����  {      9  9~�5
� �     �l�         ��t                                                                                                                                                                     c	`� 7 (    t Z� :?�          �!                                                                                                                                                                                                                                                                                                      �����                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                      �������                      �              	�          , ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$SBR2 1������ T0 �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                              � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � �                                                                                                                                                                                                                                                                                                           � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������ � ������������������������������������������������������������������������������������������������������������������������������������������������������