A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �FSAC_LST_T   8 $CLNT_NAME !$IP_ADDRESS $ACCESS_LVL  $APPS  X�$$CLASS  ������       �$FSAC_DEF_LV  ����   ������$FSAC_ENABLE         �    �$FSAC_LIST 1 ������  @!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �!�                                  �                         �