��   ?�A��*SYST�EM*��V8.2�306 4/2�
 014 A �
  ���M�N_MCR_TA�BLE   �� $MACRO�_NAME �%$PROG@E�PT_INDEX�  $OPE�N_IDaASSIGN_TYPD � qk$MO�N_NO}PRE�V_SUBy a �$USER_WO�RK���_L� M�S�*RTN � ,&SOP_�T  � �$�EMGO���RESET�MsOT|�HOLl���12�ST{AR PDI8GU9GAGBGC��TPDS�RELt�&U� �� �EST���/SFSP�C��`�C�C�NB�B�S)*$8*$3%)T ''5%)6%)7%)|S�PNSTRz�"D�  �$$C�Lr   ��i��!�����:�LDUIMT  ��������$MAXDRI�� ���%
�$.1� �% �� d%Ope�n hand 1�����%ZG_M�ENUEC?��_�x3�!(�X! %?Close3?F=p�?�?���"  �!��#S0CUST_MN �?I:�6&Oq:��6*60 ;�8d 23OO�oO8O�3(�� UB�9eO�?�O�?�3�1~�3Relax�O��OK_]_�9�6  __�_H_�_�=�"�1�_0�_�_o�_ �_Vo I:No�o�7�3Fo�ojo �o�o�o�o'�oK�o �0�Tf�� ����G��W�}� ,�>���b�׏����� ��
�C���y�(��� L�^����П	���ʟ ?��c��$�^���Z� ϯ~������)�د� $�q� ���D�V�˿z� ۿϰ�¿7��[�
� ϑ�@ώ���vψ��� ��!�����/�i�Tߍ� <�N���r��ߖߨ��� /���S����8�� \�n���������� O���_���4�F���j� ��������K�� �0�Tf�� ���G�k ,f�b���/ �1/��,/y/(/�/ L/^/�/�/�/	?�/�/ ??�/c??$?�?H?�? �?~?�?O�?)O�?�? 7OqO\O�ODOVO�OzO �O�O�O�O7_�O[_
_ _�_@_�_d_v_�_�_ �_!o�_�_Woogo�o <oNo�oro�o�o�o �oS�8� \n������ O��s�"�4�n���j� ߏ�����ď9���� 4���0���T�f�۟�� ����ҟG���k�� ,���P���ׯ����� ��1���?�y�d��� L�^�ӿ��������� ?��c��$ϙ�HϽ� l�~ϸ�ߴ�)����� _��oߕ�D�V���z� �ߞ߰�%���"�[�
� ��@��d�v����� ��!�����W��{�*� <�v���r������� ��A��<�8� \n����� O�s"4�X� ���/�9/�� G/�/l/�/T/f/�/�/ �/�/�/�/G?�/k?? ,?�?P?�?t?�?�?O �?1O�?�?gOOwO�O LO^O�O�O�O�O�O-_ �O*_c__$_�_H_�_ l_~_�_o�_)o�_�_ _oo�o2oDo~o�ozo �o�o�o%�oI�o
 D�@�dv�� �!���W��{�*� <���`���珖���� ̏A����O���t��� \�n�㟒����ȟ� O���s�"�4���X�ͯ |���ȯ�į9���� o�����T�f�ۿ�� ������5��2�k�� ,ϡ�P���tφ�������1�����
Send Event7���SENDEV�NTs��>K�� %	_�Data<��z�DATA�ߡ��=��%_�Sys�Var��|�SYS�V;��?�%G�et��<�GET���d�@w�%Re�quest Me�nu���REQMENU��۹��"� c�߇�B��Ͻ�l��� ������)��M�� �2��hz�� ��I�F. @�d����!/ /E/�/{/*/�/N/ `/�/�/�/?�/�/A? �/e??&?`?�?\?�? �?�?O�?O=O�?�? sO"O�OFOXO�O|O�O _�O�O9_�O]___ k_�_�_�_x_�_�_�_ #o�_�_okoo�o>o Po�oto�o�o�o�o1 �oU�:�� p������Q�  �N���6�H���l�� �����)��M���� ��2���V�h���� �ԟI���m��.� h���d�ٯ������� �E����{�*���N� `�տ��ҿϺ�̿A� �e��&�sϭϘ��� �ϒ�߶�+�����&��s�"ߗ�F�X��$M�ACRO_MAX��������Ж��SOPE�NBL �������y�T�T�#������PDIMSK����� �;�SU�E�W�TPDSBEOX  �S�U���߿�P�����