��   �A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG ��DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST���DwNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��,�* D� $PRIMA�R_IG !$ALTERN1�<WAIT_TI|A ��<�FT�� @� LOG�_8	�CMO>�$DNLD_FI�:�SUBDIR�CAP� W����8 . 4� H��ADDRTY�P�H NGTH�����z +L�S�&$RO�BOT2PEER�2� MASK4M�RU~OMGDE�V�W��RC�M�  $xZ ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALARl!B��TP�3�V8 S���$VAR9M� ON
6��
6APPL
6PA� 5B N	7POR��#_�!>�"ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9z!�800CH�- Y�4MAX?T��RDM*� �$DIS� *8/�SMB�	"�wBCA�$WI�2AIN4EXsPS�!�PAR��F�0BCL�
� <(C�0�SP�TMOU�4� WR8�_HuF \0@o l5��!�"�%�7X�ECC�%H� VR�0UP� �_DLV�vE(��SNo3 ��O�BX_S@~#Z_�INDE
B�QOFYF� ~UR�YD��4KT�  � t �!&PMO�N��SD��RHOU�#END�X�Q�V<�Q�VLOCA� Y�$N�0H_HE~��TCPI"�/ 3 $ARPhz&�1F�W_\ d�I!F�P;FA~qLk01#�HO_� oINFO7cEL	%G P K  !�k0WO�@ $oACCE� LVt�K�2H#ICE�>�` ��$�c# O���q��
���
�$'0 uW
���F�����ItDu�$� 2,{� ��r|} ]p�� ,}��!q����r%r,z����0�AtDq�s`_.  ,{�Krr� ��������̏ޏ�����&�8��t� _FL�TR  v4s U���������{�nx,}2�{ZbSH�w@D 1,y G P��Atџ ���2���V��z�=� ��a���ԯ������� ߯@��d�'�9���]� ����⿥��ɿۿ<� ��`�#τ�GϨ�kϡ� �������&���J�� V�1�ߤ�g��ߋ��� �����4���	�j�-� ��Q��u������ ��0���T��x�;�q�������������wz _�LI� 1]�x!1.10����0�1A��255.�y8���Iu/2 6H� \n���3�H%���
�4&H�L^p��5�H �����6/H� </0N/`/r/L�RCj`�p�p!Pp%�ː�v�� Q� ���.< (?]?o?B?�?�?�?�?�?�?��P�?O/OAO  OeOwO�O�OZO�O�O�O�.�O��Lu-_\�_�Or_�_�_�_��}�iRConnect: irc�T�//alerts �_�_oo%o�Ul_Qo@couo�o�o�o����W  �"<��d� �DM%s�~�$SMB 	���@o�/C�v�`_CL�NT 2
�� 4#T-�\�� �����3��$� i�H�����~�ÏՏ�����NM���n%�L�T��:�{��@j�����ǟ\�aN��1�m%17�2.20� 4�3�ӟ(v������8���#�UST�OM �m3����0 ���$TCWPIP�b�mX\5 TEL�e�1�2�H!TP�!�#{rj3_�tpdן # ��!KCL�諻����)u!CRT�B�0���2�!OCONS�����Osmon���