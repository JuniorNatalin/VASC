��   ,y�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_IOC_�T   P �$OPERATI�ON  $L�_TYPBIDXFBR1H[ S2]�2R�$$CL�ASS  �������P��P��$' 2 �P @ ��U���
������������������'�����  H��H� �����H� � �� �(H(D#�		/#"�H�@���H� I�=/��O�/�O�$���$ �$$%1�!� $!,5�<95 |� �<���/�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV�hz�����_C_CCL ?��� 	�All para�m��
Base��Pos./�Speed ch�eck
�Safe� I/O con/nect�}R��`���&�8�SIK�@]��r�ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m������Oʏ܏���0�+� =�O�x�s��������� ����'PK ]o������ ��(#5Gpk }����� /� //H/C/U/g/�/�/ �/�/�/�/�/�/ ?? -???h?c?u?�?�?�? �?�?�?�?OO@O;O MO_O�O�O�O�O�O�O��Nȏ  ���O&_ O_J_\_n_�_�_�_�_ �_�_�_�_'o"o4oFo oojo|o�o�o�o�o�o �o�oGBTf ��������O��SIJ����D�m� h�z�������ԏ�� ��
��E�@�R�d��� ������՟П���� �*�<�e�`�r����� ����̯�����=� 8�J�\���������Ϳ ȿڿ���"�4�]� X�j�|ϥϠϲ����� �����5�0�B�T�}� xߊߜ�������������P_8�SF'DI1�[�2a�[�I3y�[�4��[�5��[�6��[�7��[�8 ��$��'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O0�B�OF�X�O`�yCx�yC��yC�� yC��yC��yC��yC� BO3_E_n_i_{_�_�_ �_�_�_�_�_ooFo AoSoeo�o�o�o�o�o �o�o�o+=f as������ ���>�9�K�]��� ������Ώɏۏ�� �#�5�^�Y�k�}��� ����ş�����6�P1�C�NOA�SE�wB�VOFFP�FE�NCE��EXE�MG��b�ۣNT{ED�OP̯���AUTO���TO=��OݡMCyC^���CSBPv��y�dOw@A��� �����ճʯޠ��D{ISt�C_��"��_B�5�[� 