A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DMR_GRP_T  � $MASTER_DONE  $OT_MINUS   	$OT_PLUS   	$MASTER_COUN   	$REF_DONE  $REF_POS   	$REF_COUNT   	$BCKLSH_SIGN   	$EACHMST_DON   	$SPC_COUNT   	$SPC_MOVE   	$ADAPT_INER   	$ADAPT_FRIC   	$ADAPT_COL_P   	$ADAPT_COL_M   	$ADAPT_GRAV   	$SPC_ST_HIST   	$DSP_ST_HIST   	$SHIFT_ERROR  $SPC_CNT_HIS   	$MCH_PLS_HIS   	$ARM_PARAM   d$MASTER_ANG  $DSP_ST_HIS2   	$CLDET_CNT   	$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$GRAV_MAST   BL�FMS_GRP_T t *$REM_LIFE   	$NT_LIFE   	$T_LIFE   	$CLDET_ANG   	$CLDET_DSTB   	$NT_LIFE_0   	$T_LIFE_TEMP   	$REM_LIFE_0   	$GRP_CL_TIME  $PCCOMER_CNT   	$FB_COMP_CNT   	$CMAL_DETECT   	$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $DTY_STR_T  $DTY_END_T  $CLDET_CNT   	$CLACT1   $CLACT2   $CLACT3   $CLACT4   $CLACT5   $CLACT6   $CL_OVR   $CLOMEGA1   $CLOMEGA2   $CLOMEGA3   $CLOMEGA4   $CLOMEGA5   $CLOMEGA6   $CL_FRMZ   $CLDEPT_IDX   $CLCURLINE   $CLDEST1   $CLDEST2   $CLDEST3   $CLDEST4   $CLDEST5   $CLDEST6   $CLNAME ?( �PLCL_GRP_T  � 	$CALIB_STAT  $TRQ_MGN   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	P�VCAX_REFA_T  @ $REF_FACTORY  $NUM_SET  $MAST_TO_REF  $PRE_MST2REF   ��VCAX_REFD_T  , $COMMENT $REF_UPDATE  $REF_AXIS 2 	$�VCAX_REFS_T  8 $STEP_MS_ENB  $NUM_SET  $STEP_DATA  $PRE_STEP  �VCAX_REFM_T   $IS_SET  $MASTER_COUN  �VCAX_REFG_T  0 $REF_DATA 2 
$REF_STEP 2 	$PRE_MASTER 2 	�$$CLASS  ������       �$DMR_GRP 1 ������      	                                      	                                      	  1 Å�����ۢ���$ to                 	                                      	                                      	                                    	                                	  �m�HSW F�"������޽�             	                                      	                    	                    	                    	                    	 �� �:����       	   �          	 B  B   B  B                   	  i4EKt ��6I�v�R j�             	  W��  �S�۷�x� r�             d                                                                                 =L��                                    ?�                              @�                                                                                                                                                                                                                                                           	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 �����$FMS_GRP 1������  	 J���H$��F�4�J�ԓJ)0\OT��             	 M��~PI��QܼKk�K��K�7             	 B�  B�  B�  B�  B�  B�               	 BD��B&D��		�B�@��@�v��             	                                      	 N7�(P���Q��}K�ٿLLWx             	 B�vB�vB�vB�vB�vB�v             	 J��H$��F�d�J���J)0�OT��            X�Y� 	                                    	                                     	                                                                XU[
XUe:XZ&hXd�9Xh�lXh�&X�9�X�E�X���XÎ4XÎVXÎ\X�+�X�+�X�Y�XRk�XS~bXS�XTRXT�fX�(�X�)@ 	    c       '                         ��@ �� �5 �������衡 �	a ��u ����Q��-�.Y�/��,i ��< �� ��� �� �a �
x  �+H
�+=��+MG�+Y��������}�+?s�+A��+L�q�(�q�Z�q�i�q�0�q��+`U�+O!�+?$�+U��+6q�+G|   )�� )�� )�� )�� ��� �1� )� )�� )� �T� �Q# �N �,� �]� )�� )� )�� )�� )�G )�	  ���� ����iV	��P���������[5�\��\��DG�\{���7��������
  ��A��1��5��Jg�a���/����-���CM��@��R���R�l�R�g�R�~�R����K��4���8��4;��0���0  ���b�������K���x�)8�7!����+����������!���*��,���>���++���b���A������u�������     d   d   d   d      d   d   d   d   d   d   d   d   d   d   d   d   d   d   d  ���x�������0����   �  ����J�������������������    �������*��������������N����  ����������g���   G  	?�����������   ��������      B���V����������*�������[  ������������������  n����������������   ���������������*�����������'�������~  ��������������������  �����������������      ��������������������������������  ����������������������������������������          ����������������������������     S   P   b         V��������   =   <����      `   V   ]   V����   �   H   �    .  .  .  .   e   e  .  .  .   e   e   e   e   e  .  .  .  .  .  .                                                            ~                                     F                                               ?[c?[��?[�&?[�S��࿿�1$?[�E?[`�?[���h�)�iU��iU��h�-�h�v?[�S?[Ǧ?[��?[�\?[��?[�  ?:y,?9�?9�M?9�0>���>�l�?9!�?:v=?9
r?�H?�?�?�G?�-?9�0?9�?9�f?8Y�?9�?9�  ��ʾޟ�����"7������XS����}�͝B���|���|�͝9�͜���fo��ľ�۾ޟ�]  ?�ST?���?��"?��2�c�/>��?��?�S�?��?t�?t�?t�?t�?t�?��2?�W?��^?��F?���?��  ����������U���y��֌���>���S���迫Я�2�n�2��2��2�n�2�l���x��ִ��� ���A��ҽ���  ���u���Q���v�������������������ݮ���p�ÁM�ÁM���m���G������R������o���Q���.  ,($UP003                                     ($UP003                                     ($UP003                                     ($UP003                                     ($MAKRO080                                  ($UP001                                     ($UP003                                     ($UP003                                     ($UP003                                     ($MAKRO080                                  ($MAKRO080                                  ($MAKRO080                                  ($UP001                                     ($UP001...........................0020      ($UP003                                     ($UP003                                     ($UP003                                     ($UP003                                     ($UP003                                     ($UP003                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      �$PLCL_GRP 1������� D    	 ?�  ?�  ?�  ?�  ?�6?,E?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$VCAX_REF_GR 2������ t 
 �REFERENCE 1        	                                                                                                                                                 REFERENCE 2        	                                                                                                                                                 REFERENCE 3        	                                                                                                                                                 REFERENCE 4        	                                                                                                                                                 REFERENCE 5        	                                                                                                                                                 REFERENCE 6        	                                                                                                                                                 REFERENCE 7        	                                                                                                                                                 REFERENCE 8        	                                                                                                                                                 REFERENCE 9        	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE2_1       	                                                                                                                                                 REFERENCE2_2       	                                                                                                                                                 REFERENCE2_3       	                                                                                                                                                 REFERENCE2_4       	                                                                                                                                                 REFERENCE2_5       	                                                                                                                                                 REFERENCE2_6       	                                                                                                                                                 REFERENCE2_7       	                                                                                                                                                 REFERENCE2_8       	                                                                                                                                                 REFERENCE2_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE3_1       	                                                                                                                                                 REFERENCE3_2       	                                                                                                                                                 REFERENCE3_3       	                                                                                                                                                 REFERENCE3_4       	                                                                                                                                                 REFERENCE3_5       	                                                                                                                                                 REFERENCE3_6       	                                                                                                                                                 REFERENCE3_7       	                                                                                                                                                 REFERENCE3_8       	                                                                                                                                                 REFERENCE3_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE4_1       	                                                                                                                                                 REFERENCE4_2       	                                                                                                                                                 REFERENCE4_3       	                                                                                                                                                 REFERENCE4_4       	                                                                                                                                                 REFERENCE4_5       	                                                                                                                                                 REFERENCE4_6       	                                                                                                                                                 REFERENCE4_7       	                                                                                                                                                 REFERENCE4_8       	                                                                                                                                                 REFERENCE4_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                         