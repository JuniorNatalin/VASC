��   �P�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�RYRUN_T   � $'�ENB 4 NU�M_PORTA �ESU@$ST�ATE P TC�OL_��PMPM�CmGRP_MA�SKZE� OTI�ONNLOG_IgNFONiAVc�FLTR_EMP�TYd $PRO�D__ L �ESTOP_DSBLA�POW_RECO�VAOPR�SA�W_� G %�$INIT	RE�SUME_TYP�ENx&J_ � 4 $($FST_IDX��P_ICIװ�MIX_BG-yA
_NAMc �MODc_US�d�IFY_TIv� wMKR-�  $LI�Nc   �_7SIZc?\x� �k. , $?USE_FL4 ���&i*SIM�A�Q#QB6'S�CAN�AXS+I�NS*I��_COU�NrRO��_!_?TMR_VA�g�h>�i)  �'` ��R��!�+�WAR�$}H��!{#NPCH���$$CLASS  ���01��5��5�6/ 05_5�����Ec����\1l510�71p5��%VAGh���<�0TPd�?��A5I2L;�c ��"��	A$*��Y4d��Y3	A�[2)Y3�Y4-D U&H��&G\0$pAhF	~ChF�ChF�ÞChF�n@�fH�T�ChF�n@�fH�n@E�&GAA4B�D!z0�8�H`0Q�Fhz0iR�Hl.S�Fyz0��HU�z0��H�z0��H5�z0�&G~SxV	~P�HU@�QxVa@�2vX9~P;vXA�~PPvXa~PxvX�T�SxV�~P�vX�c�xV�~P�vX�@�vX�>cxV�~P�@xV)�^c(E\0Phf�=@+fhC�chfHH# �5maL�chfQ# YqfhAP{fh��c"hf�# QPhf��chfbaPqPhf�@�fh��# Eh�>s(E��@PqHvP3Fx7�nsHv�0�qHv�PsFxw�sHv��sHv!`��Fx1p�&GH�@�q�v �s�v1�pD�P�vV�p�P�vv�p����=AD��G&�M����U=AAP z&�T^�)�����&��~�T)��q�&����&�����&�ae=A�P��eU=A�A�&����,�@(� ��P ����P ���J.���@�P@����PP���` $U��en���u �UP��U������ �&�#
n@�P(���DB
���z0��?���������6W?05�V1 F�OLGE��U��U  0h�MA�KROa�SUCyH�eh�BIN����D�o { 2}L; 4%|��SP��ׯ���J�{�IƦ�U
�  �</t�̠eu>� ' h=eq%�}1Ʀ4A���5-��Y�;2L����="k���6����\�uu�  am`u���UB����"� ����L?������X�P$�"�X �01�\0�0tq*� _t
 Nq��P����F������ �1�C�U�g�yߋߝߐ�>i5}1��s����B�qu) H��I�qs��Zr��\t{tq�иttt}1 �'�9�K�]�o���������7� �2t� � ����&�8�J�\�n� ��������������i7 �,>Pbt� �������� (:L^p��� ���� /$/6/ H/Z/l/~/�/�/�/�/ �/�/�///2?D?V? h?z?�?�?�?�?�?�? �?
O?.O@OROdOvO �O�O�O�O�O�O�O_ _#O<_N_`_r_�_�_ �_�_�_�_�_oo_ 1_Jo\ono�o�o�o�o �o�o�o�o"-oF Xj|����� ����0�;T�f� x���������ҏ��� ��,�7�I�b�t��� ������Ο����� (�:�E�^�p������� ��ʯܯ� ��$�6� H�S�l�~�������ƿ ؿ���� �2�D�O� a�zόϞϰ������� ��
��.�@�R�]�v� �ߚ߬߾�������� �*�<�N�`�k߄�� �����������&� 8�J�\�g�y������ ��������"4F Xju������ ��0BTf x������� //,/>/P/b/t/ ��/�/�/�/�/?? (?:?L?^?p?�?�/�? �?�?�?�? OO$O6O HOZOlO~O�O�?�O�O �O�O�O_ _2_D_V_ h_z_�_�O�O�_�_�_ �_
oo.o@oRodovo �o�o�_�o�o�o�o *<N`r�� ��o�����&� 8�J�\�n�������� �ڏ����"�4�F� X�j�|���������֟ �����0�B�T�f� x���������˟��� ��,�>�P�b�t��� ������ǯٯ��� (�:�L�^�pςϔϦ������ջ ds_
 q����t���"�4�F� X�j�|ߎߠ߲����� ٿ����0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ������$6 HZl~���� ��� /2/D/V/ h/z/�/�/�/�/�/�/ �//?.?@?R?d?v? �?�?�?�?�?�?�?O ?*O<ONO`OrO�O�O �O�O�O�O�O_OO 8_J_\_n_�_�_�_�_ �_�_�_�_o_4oFo Xojo|o�o�o�o�o�o �o�o)oBTf x������� ��%7P�b�t��� ������Ώ����� (�3�L�^�p������� ��ʟܟ� ��$�6� A�Z�l�~�������Ư د���� �2�=�O� h�z�������¿Կ� ��
��.�@�K�d�v� �ϚϬϾ�������� �*�<�N�Y�r߄ߖ� �ߺ���������&� 8�J�U�g߀���� ���������"�4�F� X�c�|����������� ����0BTf q�������� ,>Pbm ������// (/:/L/^/p/{�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�/�?�?�? �?�?�?O O2ODOVO hOzO�?�?�O�O�O�O �O
__._@_R_d_v_ �_�O�_�_�_�_�_o o*o<oNo`oro�o�o �_�o�o�o�o& 8J\n���o�o �����"�4�F� X�j�|������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ǟ���� (�:�L�^�p������� ��ïܿ� ��$�6� H�Z�l�~ϐϢϴ��� ѿ����� �2�D�V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����������& 8J\n���� ������"4F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ /?,?>?P?b?t?�? �?�?�?�?�?�?�/? (O:OLO^OpO�O�O�O �O�O�O�O _O$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o_2oDoVo hozo�o�o�o�o�o�o �o
o'o@Rdv �������� �#<�N�`�r����� ����̏ޏ����&� 1�J�\�n��������� ȟڟ����"�-�?� X�j�|�������į֯ �����0�;�T�f� x���������ҿ��� ��,�>�I�b�tφ� �Ϫϼ��������� (�:�E�W�p߂ߔߦ� �������� ��$�6� H�S�l�~������ ������� �2�D�V� a�z������������� ��
.@R]�o� ������� *<N`k�� �����//&/ 8/J/\/n/y�/�/�/ �/�/�/�/?"?4?F? X?j?u/�/�?�?�?�? �?�?OO0OBOTOfO xO�?�O�O�O�O�O�O __,_>_P_b_t_�_ �O�_�_�_�_�_oo (o:oLo^opo�o�_�_ �o�o�o�o $6 HZl~��o�� ���� �2�D�V� h�z������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ��ڿ����"�4�F� X�j�|ώϠϲϽ�Ͽ ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p��������������� _ds
�qu����q����qs�s����tr� t�� q �t��CUgy����������`V��J L K �Mquqs)�Arskq) �t!;'�tt1K ]o������\���ads���,[�r8tB, � u(H""I Z  \9J/\/n/ �/�/�/�/�/�/�/�� ?"?4?F?X?j?|?�? �?�?�?�?�?�??O 0OBOTOfOxO�O�O�O �O�O�O�OO_,_>_ P_b_t_�_�_�_�_�_ �_�_o_(o:oLo^o po�o�o�o�o�o�o�o  o6HZl~ �������� 2�D�V�h�z����� ��ԏ���
��'� @�R�d�v��������� П�����*�5�N� `�r���������̯ޯ ���&�1�J�\�n� ��������ȿڿ��� �"�4�?�X�j�|ώ� �ϲ����������� 0�B�M�f�xߊߜ߮� ����������,�>� I�b�t������� ������(�:�L�W� p���������������  $6HZe�~ �������  2DVaz�� �����
//./ @/R/d/o�/�/�/�/ �/�/�/??*?<?N? `?r?}/�?�?�?�?�? �?OO&O8OJO\OnO y?�O�O�O�O�O�O�O _"_4_F_X_j_|_�O �_�_�_�_�_�_oo 0oBoTofoxo�o�_�o �o�o�o�o,> Pbt��o��� ����(�:�L�^� p��������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ�ſ�� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ���(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�?  ?2?D?V?h?z?�?�? �?�?�?�?�/
OO.O @OROdOvO�O�O�O�O �O�O�O�?_*_<_N_ `_r_�_�_�_�_�_�_ �_o_&o8oJo\ono �o�o�o�o�o�o�o�o 	o"4FXj|� ������� 0�B�T�f�x������� ��ҏ�����%�>� P�b�t���������Ο �����!�:�L�^� p���������ʯܯ�  ��$�/�H�Z�l�~� ������ƿؿ����  �2�=�V�h�zόϞ� ����������
��.� 9�R�d�v߈ߚ߬߾� ��������*�<�G� `�r��������� ����&�8�J�U�n� ���������������� "4FQ�j|� ������ 0BT_x��� ����//,/>/ P/b/m�/�/�/�/�/ �/�/??(?:?L?^? i/�?�?�?�?�?�?�?  OO$O6OHOZOlOw? �O�O�O�O�O�O�O_  _2_D_V_h_z_�O�_ �_�_�_�_�_
oo.o @oRodovo�_�o�o�o �o�o�o*<N `r��o���� ���&�8�J�\�n� �������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϱ�������  ��$�6�H�Z�l�~� �ߢߴ߿��������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/��/?? 0?B?T?f?x?�?�?�? �?�?�?�/OO,O>O PObOtO�O�O�O�O�O �O�O�?_(_:_L_^_ p_�_�_�_�_�_�_�_ �Oo$o6oHoZolo~o �o�o�o�o�o�o�oo  2DVhz�� �����
�.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ����8�J�\�n� ��������ȯگ��� �"�-�F�X�j�|��� ����Ŀֿ����� )�B�T�f�xϊϜϮ� ����������,�7� P�b�t߆ߘߪ߼��� ������(�:�E�^� p�����������  ��$�6�A�Z�l�~� ��������������  2DO�hz�� �����
. @R]v���� ���//*/</N/ Yr/�/�/�/�/�/�/ �/??&?8?J?\?g/ �?�?�?�?�?�?�?�? O"O4OFOXOjOu?�O �O�O�O�O�O�O__ 0_B_T_f_qO�_�_�_ �_�_�_�_oo,o>o Poboto_�o�o�o�o �o�o(:L^ p��o�����  ��$�6�H�Z�l�~� �����Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤϯ��������� �"�4�F�X�j�|ߎ� �߲߽��������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p��������  $6HZl~ �������/  /2/D/V/h/z/�/�/ �/�/�/��/
??.? @?R?d?v?�?�?�?�? �?�?�/OO*O<ONO `OrO�O�O�O�O�O�O �?__&_8_J_\_n_ �_�_�_�_�_�_�_�O o"o4oFoXojo|o�o �o�o�o�o�o�oo 0BTfx��� �����,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ���6�H�Z�l�~� ������Ưد���� �2�D�V�h�z����� ��¿Կ���
��'� @�R�d�vψϚϬϾ�@��������*� 