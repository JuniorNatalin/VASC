��   t��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���U�I_CONFIG�_T  d �9$NUM_MENUS  9�* NECTCRE�COVER>CCOLOR_CRR�:EXTSTAT���$TOP>_�IDXCMEM_�LIMIR$D�BGLVL�PO�PUP_MASK��zA  $DUMMY54��ODE�
5CFO�CA �6CPS�)C��g HA�N� � TIME�OU�PIPES�IZE � MW�IN�PANEM;AP�  � � �FAVB ?� 
w$HL�_DIQ�?� qELEM�Z�UR� l� S|s�$HMI��RO+\W AD�ONLY� �T�OUCH�PRO�OMMO#?$��ALAR< �F�ILVEW�	E�NB=%%fC �1"USER:)FC[TN:)WI�� I* _ED�l"V!�_TITL� ~1"COORDF<#/LOCK6%�$F%|�!b"EBFOR�? �"e&
�"�%�!�BA�!j ?�"B�G�%$PM�X�_PKT�"IHE�LP� MER�B�LNK$=ENAB��!? SIPMAN�UA�-4"="�B�EEY?$�=&q!E�Dy#X&UST�OM0 t �$} RT_SPI�D��4C�4*PA�G� ?^DEV�ICE�9SCREVuEF���7N��@$FLAG�@�%�1  h �	$PWD_ACGCES� E �8��TC�!�%)$L�ABE� 	$T�z j4@q!�D�	��&USRVI| 1  < ` �B��APR�I�m� U1�@T�RIP�"m�$$�CLA?@ �����A��R��R��$'2 ~����R�	 ,R��?���/Q=Q(8R3T.Q��
��)P�  1T<w_��
 ���A�_@�_�_�_�_�_o �_ *o<oNo`oro�oo�o �o�o�o�o�o&8�J\n���(/�SOFTP�0/G�ENLINK?c�urrent=m�enupage,935,1��� ��!:�L�^�p��� ��#���ʏ܏� �� ��6�H�Z�l�~����� 1�Ɵ؟���� ����D�V�h�z�������� TPTX�����:�ٯ�� s� Ƿ���$/s�oftpart/�genlink?�help=/mdw/tp�q.dg�� F�X�j�|�5�&�#�pwd2�ɿۿ��� 4�#�5�G�Y�k�}�� �ϳ��������ϊϜπ1�C�U�g�yߋ�aT���AoP��QR�� ($ ����������(����A2QN�PSHr_PS���^�
q��2Q����RQ  ���ʡ��	�������L�L�Y��S�2 1�E=PR_ \ }�mPREG V�ED��6�H�wh�olemod.h�tm\�singl�m�doub���trip��brows����I� ������3EWi�{�3�W�i�dev.sr�l���	1�	t ��	� �o��]���8��(/� �@@/ R/d/v/�/�/�/�/�/�/�& @</?#?�/ G?Y?k?:6+�#//�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O��O�O#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo 5/�o�o�o�o�o�o  2D??hzI[ ��y?�?qo
��� )�R�M�_�q������� ���ݏ��*�%�7� _W�Q��������ǟ ٟ����!�3�E�W� i�{�������ï�o�� �"�4�F�X�j�|��� ���Ŀֿ������ ��ͯf�a�sυϮ� �ϻ���������>� 9�K�]߆߁ߓ�a��� ���������#�5�G� Y�k�}�������� �������Z�l�~� ����������������  2hz1�C� )�����
 )RM_q��� ������/	/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?I��?�?�?�?�? O"O4OFOXOS|O�O�]OoO�O�O�J�$U�I_TOPMEN�U 1�@Q�R 
X�Q�1)*def�ault�?�=	�*level0 *HP 8_& o_�_m_Rtpio�[23](tpst[1�X�_�_�_�BVX_�_!$
h58e01.gifo~(	menu5Bi9`da13BjcbAjad14ikPoa���o�o �o $6�2�o_�q����Htp�rim=dapag�e,1422,1 ����/�A�Le�@w���������N��vclass,5ȏ@���!�3�E�P�܌13L���������ʟQ��|53���P*�<�N�Q��|8�� ��������ѯP���� �+�=�O��9PQ _��B]y�aw��oÿƹVty�]�_�Qmf�[0�_��	�c[g164�W>�59�X a�oٿ{�]h2�ogm ��}j�osgAk���cg� y�F�X�j�|ߎ�寲� ����������0�B�@T�f�x���ۍ2�� �����������O� a�s�����&�8�p���@���� ۟�14�@^p���%��s?ainedi����%�wintp�p0bt�� ��6Qr���fo ��//0/B/T/f/x/ �/ o�/�/�/�/�/? ?,?>?c?�o�?�?�? �?�?�? �OO)O;O MO_O�?�O�O�O�O�O �O�O~O_%_7_I_[_ m_�O�_�_�_�_�_�_ z_o!o3oEoWoio{o 
o�o�o�o�o�o�o�o /ASew��������� o�0������⯿]?o���s󽌏������u ��d�f���&�4�����B�h��ό�6��u7 ���0����'�9� �]�o���������F� ۯ����#�5�G�64�1C��������� ɿԯ����#�5�G� ֿk�}Ϗϡϳ����� 2�����1�C�U�����6\ߑߣߵ�����4Ӝ74��'�9� K�]�������/z� ���������"�G�F� ��R�|����������� ����p?1CUgy �Vϯ����	 �?Qcu�� (����//� ;/M/_/q/�/�/�/6/ �/�/�/??%?�/I? [?m??�?�?2?�?�? �?�?O!O3O�?WOiO {O�O�O�Ol�~��O�� l�
_._@_R_w_v_ �_�__�_�_�_oo o*o<oNo�o�o�o �o�o�o�oHO'9 K]o�o���� ��|�#�5�G�Y� k�}������ŏ׏� �����1�C�U�g�y� �������ӟ���	� ��-�?�Q�c�u���� ����ϯ����O�O ;��O�_^op������� ��ʿܿ�\���7�6� H�Z�l�~ϐϢ�po�� �����!�3�Eߜ�i� {ߍߟ߱���R����� ��/�A�S���w�� ������`����� +�=�O���s������� ������n�'9 K]������� �j�#5GY k&����ϲ��� ��//0/B/�b/ `/�/�/�/�/�/�/�/ ?��??Q?c?u?�?�? ��?�?�?�?OO�? ;OMO_OqO�O�O�O6O �O�O�O__%_�OI_ [_m__�_�_2_�_�_ �_�_o!o3o�_Woio {o�o�o�o@o�o�o�o /�oSew� ���z���? ?*�<�N�`�r����� �����ޏ����&� K�J�\�*?������ɟ ۟�D�#�5�G�Y� k�}������ůׯ� �����1�C�U�g�y� �������ӿ���	� ��-�?�Q�c�uχ�� �Ͻ�������ߔ�)� ;�M�_�q߃ߕ�$߹߀���������w�t�*default��w�*leve�l8ˏi�{��7� �tpst[1�]����y��tpio[23������u��n��6�H�	m�enu7.gif�I�
h�13m�z�5Ђ�g��e�4��u6 m�����%7I ��m����V ��!3EW��prim=h�p�age,74,1�\�������pclass,13�/(/:/L/^/��5d/�/�/�/�/�/���/?.?@?R?d?gy18��?�? �?�?�?�/�6�?%O�7OIO[OmOL��$U�I_USERVI�EW 1�q�q�R 
���tON�O�OF�m �O__%_7_I_�Om_ _�_�_�_X_�_�_�_ o!o�O.o@oRo�_�o �o�o�o�oxo�o /AS�ow��� �jo���b+�=� O�a�s��������͏ ߏ����'�9�K���*zoom^�ZOOM]���� ԟ���
���.�@�R� d�v��������Я����*maxr�es��MAXRES������\�n��� ����G�ȿڿ���� ��4�F�X�j�|�'��� �ϭ��������0� B���f�xߊߜ߮�Q� ����������'�=� K�߆������q� ����(�:�L���p� ��������c������� [�$6HZl� ����{�  2D��Ucu�� ����
/�./@/ R/d/v//�/�/�/�/ �/��/??�/N?`? r?�?�?9?�?�?�?�? OO�?8OJO\OnO�O #A