A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DCSS_CPC_T   � $COMMENT $ENABLE  $MODE  $GRP_NUM  $MODEL_NUM   $UFRM_NUM  $NUM_VTX  $X   $Y   $Z1  $Z2  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD  �DCSS_CSC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $TCP  $UFRM_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  �DCSS_GRP_T  � $TCPCHG_SIZE  $APSPD_MODE  $ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $APSPD_JMODE   	$ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$TCP_SEL  �DCSS_GSTAT_T  D $FP_BASE $LINK_BASE ! 	$LINK_BASE_V ! 	$LINK_BASE_H ! 	 !�DCSS_JPC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $UPR_LIM  $LWR_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD   �DCSS_JSC_T  | 
$COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  ��DCSS_ELEM_T  T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    %��DCSS_MODEL_T   $COMMENT $ELEM 2 
�DCSS_PSTAT_T  � 	$STATUS_CPC    $STATUS_CSC   $STATUS_JPC   ($STATUS_JSC   ($USER_MODEL   $ROBOT_MODEL   $USER_ELEM   $ROBOT_ELEM   $CUR_TCP   $�DCSS_SETUP_T 	 l $DISP_MGN  $INP_ASSIST  $TOOLCHG_ENB  $DO_TYP  $DO_IDX  $DO_MGN  $CALMD_ENB  $CALMD_STAT  ��DCSS_T1SC_T 
  $ENABLE  $SPD_LIM  �DCSS_TCP_T  l $COMMENT $UTOOL_NUM  $MODEL_NUM  $VRFYIO_TYP  $VRFYIO_IDX  $X  $Y  $Z  $W  $P  $R  ��DCSS_SPH_T  ( $SIZE  $DATA1  $DATA2  $DATA3  �DCSS_BOX_T  8 $SIZE1  $SIZE2  $SIZE3  $X  $Y  $Z  $R  ��DCSS_TUIRO_T  , $TYPE  $SPHERE 2 $BOX $BOX_S 2 ��DCSS_TUIZN_T  0 $ENABLE  $X   $Y   $Z_UPR  $Z_LWR  �DCSS_UFRM_T  @ $COMMENT $UFRM_NUM  $X  $Y  $Z  $W  $P  $R  $�$$CLASS  ������   Q    Q�$DCSS_CPC 2 ������Q   ��                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �$DCSS_CSC 2������Q  D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_GRP 2������Q  �                         	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                         �$DCSS_GSTAT 2������Q  ,8�?L���9�>�M���/ӿic=C7�>�Qݾx���]�KD������D�D/��� 	 88�?h��`j    4r�4��8?�  ��`j�h4��ZC�bt���    ���8��!'�=�J�?|c�d}�>��1�G��`j�h4��ZB�-Z�S��D�Uf���8����>X`R?]��>�`b?h���x�H�>�c:����A:�����D������8���Q�>x��?]�L�H�>�cC���о�X:�e�]<���D~g���D찻���8�?H�cB>���>�X5?e�^���h��Q�>x��?]�KD~g���D찻���8�?L���9�>�M���/ӿic=C7�>�Qݾx���]�KD������D�D/���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8���������������������������������������� 	 88����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8����������������������������������������8�����������������������������������������$DCSS_JPC 2������Q ( D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_JSC 2������Q ( @BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                               =���BS HALT                                               =���BS HALT                                 	              =����                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �$DCSS_MODEL 2������Q x�                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �$DCSS_PSTAT ������Q       (  (     ����                                                                                    ������������                  �������������$DCSS_SETUP 	������QB�                B�          �$DCSS_T1SC 2
������Q      Cz      Cz      Cz      Cz      Cz      Cz      Cz      Cz  �$DCSS_TCP R������Q � 
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �$DCSS_TCPMAP  ������Q @                            	   
                                                                      !   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @�$DCSS_TUIRO 2������Q �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$DCSS_TUIZN 2������Q 	 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �$DCSS_UFRM R������Q � 	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      