��   v��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<�$1_8k 8��FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\9 ^75z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D��VCAX_�w A.  @ 5vFX0OR�@E ?NUM_SE238�_TO0Q�#RE_:� 2cT |+V>1 , $� �ME�vUPgDAT�wAXy_2 	�+VS5Q' 8<P��PnP;0k L\�R�PA�kQ�Q��+VM5Q  �$ISRTd 5+VG5Q { v��R2 
v�S2�T kR9�P 	��$U1SS  O����a����w�$' 1 �e� } �� 	 ����o�o�o�f|]�;�Cq�����  W��*�j�o�oA,ePz���yM}�a��|���8����?�`q+ �4���9����T� ����|�+�=�d��a�����%���CZ� ������wBgB ���`B���f��p���z3�������;�����$ �]�o~	��Q����W^p�p�
pA��d�1�C�U����=L��`���?�����@���͟ߟ ���'�9�K�]�o������� �e��̧8��쯄d  2 �� /�A�S�e�w�����������<������ 1�C�U�g�yϋϝϯ� ���`�a�o������ *�<�#�`�K߄�oߨ� ��c��ߡ����&�[� 5�G�n�k�}����� ��������"���P� b�t������������� ��(:��^p ������Eϯ� �6HZl~� ����˿�/ / 2/D/V/h/z/�/�/�/ �/�/���/��/.?? R?9?v?a?�?�?�?�? ���?�?OO<O'O�? ]OoO�O�O�O�O3O�O �O_�O_J_=�k_}_ �_�_�_�_�_�_�_o o1oCoUo|o�o�o �o�o�o�goio�o- #Tfx���� �����,�>�P� b�t���������Ώ�� ��/�(��L�7�p� W������ʟ����? �՟6�!�Z�l��O{� ������ïկQ���� 2�D�/�h�[_������ ��ѿ�����+�=� O�a�s�5�ϬϾ��� ����G���'�K�A r߄ߖߨߺ������� ���m�J�\�n�� ����������������$FMS_G�RP 1^� >��I��$Gr�D�H�eIt��I��uI4l�J�M+�P�~��PxK���J��LJ��=pJ�B�  ����B��LB!v����y�?�\����A�j�J����u��)�Q�:�BP˙K���Ke��Kw\�e���X?�X��O�Gs��H�It��#I��I5=�+�X�5��������/���N3� �U� �  4� U!}�U#!z?��C�?�Vsa��S�S�V�DU__!_&� �ËNuF�N���oQO�T��,�U!{aX뿽HX���
4�4�0��8��q� �A� ����� ����<������87s86��7�b7������t���n�;U�rB���N�,����6�7 3!��������#����: ��x0 �B� ��L�����J�-��:�Nq)�N� �{O �.^E �u� |6�ҵ�7������9o#�=�Ù������������~ ��k� ȱG ���� �����Rm�b� �a'�����{���։�BB�"�P�����M�#���� ���/���c������8�������~N�ׂ���^��Z���� �H1��n�Đ� �譻4Q����@��U�3�����"F'0C�"E����d��I����!o��.�a���I����h�NN��4����!L�Z�$��`�7���B��\~�g0��k3Fs0�v�.�x��y�������������������~BV�~A����i��J��������[%N"}�  �4
5i��7��1�9�1�?}��2�
_��_��D��_е�,@�
�#���w4�+_��  �,@>  t w ��� �+AT�5cD_��4����4�GC�z@�"4���� � ��0\���-�[C��4�D^@�B�_��_��_��  8_Э�0EV
��4�M���@e,�0��0�'8�3Q2A.@�B�
�_Б��
�_иA4�WVkC��_��_�� @���06PZ@PD��_Ъ@V�1!_�ʹ
����>,@����0� @�  ��  g)�3�%_��TfA���
�&_ОP 9
�Ս�TAW@,@����  �z�4A��?o'o1fiȳ4Yoko}o �Q�o�3
�1�8	�d�5�1�*�i�d�4!4��A�7?%�B�.*�mY�r���9��c����꿪�����P�����������)���`�?�7A?��5b��
?"��*��� ��ߏ�>�R
2����>�ھ>���[r��>��5��������%�ڐ�>��q>���>��P�>���?7���?4[>�l��˾�1���B��3ҿt����b�[��ÿC���<�s�y��A�������8x��2���nT�
~�ʿp��
=��ʦK��N�_��:�?���ʾ����QF�d?l��7���%�啤���$�b����O?�#y?�����������@׿�`ƿ���/<�>G<��3&?��<���?�?��t�"��r�W���᯿��d�W�e������e�o�e���e�%�����S�����y����]~���ƿ��8��W%ҿ��S����������bH�K?��-?�"e����?�#�����u迀�@$�{�@%��@$�@$��?�^�?jq���}�?K�
����x��:�����%	,($UP�003�o� ��1 �;�"�_�F���j�|�`����ݟğ��2.��א8��6��/�A��ϓFOLGE124g�s����������� ˯ݯ�͙��J�1�n� ��y���^�ǿ���ҿ �!��EϨVo{�f� �ϊ��Ϯ������� �A�,�e�P߉�p߂� �ߪ�������U/� A�Toe�w����߿� N���������=�O� a� ���������z��� ����9K] ����v��� �5GY}� ��r���/� 1/C/U//y/�/�/�/ n/�/�/�/	?�/-???�Q??u?�?�?�?*A� o?�?�?�?c?O.O@O ROOvO�O�O�OkO�O �O�O�O_*_<_N__ r_�_�_�_g_�_�_�_��\��1234567890o'e��o Io9omo]oyo�o�o�o �o�o�o�o!-5 G{k����� �����S�C�_� g�y���������ӏ� ����7�a���� �����ӟ���0� �T�?�x�c�u����� ү������,�#�P� �_t�������	���� o���(��L�^�p� ��AϦϸ����ϛ� � �$���H�Z�l�~�=� �ߴ����ߗ���� � ��D�V�h�z�9��� �������
����@� R�d�v�5��������� ������<N` r1����?�� 8J\n- �������/ �4/F/X/j/)/�/�/ �/�/�/�/�/?oc� 9?Q�]?M?i?q?�?�? �?�?�?�?OOO%O 7OkO[OwOO�O�O�O �O�O�O�O_C_3_O_ W_i_�_�_�_�_�_�_ �_oo'oQoAouou� ?�o�o�o�o�o�o  D/Aze�� �������@� 7�d�v��/������Џ /�􏃏�*�<�N�� r�����U���̟ޟ� ���&�8�J�	�n��� ��Q���ȯگ쯫�� "�4�F��j�|���M� ��Ŀֿ迧���0� B��f�xϊ�IϚ��� ���ϣ���,�>��� b�t߆�Eߖ߼����� ���(�:��^�p� ��A�������� � �$�6���Z�l�~�=� ������������  2)?MeoYas� ����� '[Kgo��� �����3/#/?/ G/Y/�/}/�/�/�/�/ �/�/�/?A?1?e?U?�q?y?�1�$PLC�L_GRP 1����1�� D�0�?��  �:w�'?o��9�O�:O %O^OIO�OmOO�O�O �O�O _�O�>2_�OY_ �O}_h_�_�_�_�_�_ �_�_o
oCo*o$_vo 8o�o4o�o�o�o�o	 ?*cN�n ho�|�x��)� �M�_�J���n������ˏ=�$VCAX�_REF�0 2��5 �t 
 ����ERENCE 1��׏7�I�[�m�������2�ԟ柀��
��.�@����3 ß|�������į֯�S��4k�$�6�H�Z� l�~������5�̿ ޿���&�8ϣ�� �4��zόϞϰ������ϱ�7c��.�@�R� d�v߈����8��� ��������0���9��l�~���������C�FACTORY DATA\� �'�9�K�]�o������9������������	 ��GYk
�2_����������2_ �Pbt��� �'j�?�
//./ @/R/d/'���/�/ �/�/�/�/?'���/ H?Z?l?~?�?�?�?' b�7?�?OO&O8OJO \O'
��?�O�O�O�O �O�O_'�ՇO@_R_ d_v_�_�_�_'Z�/_ �_�_oo0oBoTo�� �_�o�o�o�o�o�o�o ��/ASew@%�����3� �%�7�I�[�m���_ �t7��Ώ����� (������d�v����� ����П;����/�� 0�B�T�f�x�㟥�/? ��Ưد���� ��� ���?\�n��������� ȿ3���O��(�:� L�^�p�ۿ��'_�Ͼ� �������߃ϥ��_ T�f�xߊߜ߮���_o qo����,�>�P�b� t������������(�:�L����4 ��������������� *�p���0BTfx ��S����  2D���� ������W ��(/:/L/^/p/�/�/ �K��/�/�/?? *?<?�/�x?�?�? �?�?�?�?O?�� O 2ODOVOhOzO�O�? C��O�O�O�O_"_4_ ����j_|_�_�_�_�_ �_�_��	�o!o3oEo Woio��o�o�o�d