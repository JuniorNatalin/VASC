A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �BIN_CFG_T   X 	$ENTRIES  $Q0FP  $Q0NP  $Q1FP  $Q1NP  $Q2FP  $Q2NP  $PPPP  $CNETP   ��DHCP_CTRL_T  0 $ENABLE  $IPUSE  $RETRATE  $SETHOST  �,�DNSS_CFG_T  8 $ENABLED  $IFACE_NUM  $DBG_LEVEL  $DOM_NAME !���DNS_CFG_T  D $PRIMAR_IP !$ALTERN_IP !$RETRIES  $WAIT_TIME  $ENABLE  ��FTP_CTRL_T  @ $LOG_ENTRIES  $LOG_CMOS  $DNLD_FILTER  $SUBDIRCAPS   t�HOSTENT_T  4 $H_NAME !$H_ADDRTYPE  $H_LENGTH  $H_ADDR !��PPPCFG_LST_T  D $ROBOTIP !$PEERIP !$NETMASK !$MRU  $COMP  $DEVTYPE   J�RCMCFG_T �  $RCM_ENABLE  $QSIZE  $TIMER  $STATUS_TIME  $MAILSERV  $PLANT <$LINE <$CLUSTER <$TOADDR P$CCADDR P$FRADDR P$SUBJECT $STATUS_ENB  $ALARM_ENB  $TPLOG_ENB  $LOG_EVENTS   $VARLOG_ENB  $MOTION_ENB  $SYSTEM_ENB  $APPL_ENB  $PASS_ENB  $COMM_ENB  $PORT  $STAT_SUBJ $ALERTADDR P$ALERTURL }$STAT_ATTACH }$ERR_THROT  $USR_THROT  $SIZE_THROT  $VARCHG_TIME  $VARCHG_MAX  D�RDM_CFG_T   $DISABLE   ~(�SMB_T 	 D $ENABLE  $BCAST  $WINS_IP !$DOMAIN !$EXPSRV  $SPARE  ��SMB_CLNT_T 
 < $CACHE  $RSPTMOUT  $SETPWRD  $DOMAIN !$SPARE   �SMTP_CTRL_T  l 	$ENABLE  $SERVER %$PORT  $TIMEOUT  $CC_ADDR %$FROM_ADDR %$RT_ADDR %$POST_DLVR  $SPARE  ��SNTP_CFG_T  X $ENABLE  $SERVER %$TIME_WIN  $TZ_INDEX  $TZ_OFFSET  $CUR_OFFSET  $DST  ��SNTP_CUSTOM_  t $START_MONTH  $START_DATE  $START_HOUR  $END_MONTH  $END_DATE  $END_HOUR  $LOCAL_TIME  $NORTH_HEM  �TCPIPCFG_T  X $ARPSIZE  $HOST_IPF  $HW_MCFILTER  $DEF_INTERFA  $CLASSMASK  $SHO_NETINFO  �TEL_LST_T  P $DEV_NAME !$PASSWORD  $ACCESS_LVL  $TIMEOUT  $PORT  $DEVICEUSE   ��$$CLASS  ������   
    
�$BIN_CFG  ������
�   F                           �$DHCP_CTRL 2������
�             
               
    �$DNSS_CFG ������
�        !�                                  �$DNS_CFG ������
�!�                                  !�                                           �$DNS_LOC_DOM  ������
� �                                                                                                                                                                                                                                 �$ETH_FLTR  ������
�        �   �            �$FTP_CTRL ������
�   2            �$HOST_SHARED 1������
  P!�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  �$PPP_LIST 1������
�  x!1.1.1.10                          !1.1.1.11                          !255.255.255.0                       �      !1.1.2.10                          !1.1.2.11                          !255.255.255.0                       �      !1.1.3.10                          !1.1.3.11                          !255.255.255.0                       �      !1.1.4.10                          !1.1.4.11                          !255.255.255.0                       �      !1.1.5.10                          !1.1.5.11                          !255.255.255.0                       �      !1.1.6.10                          !1.1.6.11                          !255.255.255.0                       �      �$RCMCFG pI�pMl
       
  � Q� �                                  <�                                                              <�                                                              <�                                                              P�                                                                                  P�                                                                                  P�                                                                                  �                                                                   �                          P�                                                                                  }iRConnect: irconnect://alerts                                                                                                 }�                                                                                                                                      0    <   d�$RDM_CFG ������
�    �$SMB 	������
      !�                                  !�                                          �$SMB_CLNT 2
������
  4          !�                                                !�                                                !�                                                !�                                                !�                                                !�                                                !�                                                !�                                      �$SMTP_CTRL ������
   %�                                            %�                                      %�                                      %�                                             �$SNTP_CFG ������
�   %172.20.254.203                              ��������   �$SNTP_CUSTOM ������
�            
            �$TCPIPCFG ������
�                     �$TEL_LIST 1������   
�  H!TP                                rj3_tpd                  ����   !KCL                               �                                !CRT                               �                         ����   !CONS                              rj3_smon                 ����   