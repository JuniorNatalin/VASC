��   ɋ�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_CPC_�T   � �$COMMENT� $ENA�BLE  $�MODJGRP_�NUMKL\ � $UFRM�\] _VTX �M �   $Y��Z1K $Z2��STOP_TY}PKDSBIO��IDXKENBL?_CALMD�&}S. � 8�J\TC�u
SPD_LI_����COL�&Y0 � � !CHG�_SIZ$A�P7ECDIS � � �7�C�����Jp 	�J �� ��"��$�'"_SEs��,xSTAT/� D $FP_�BASE �$LINK`$!��j&_Vs.Hs#�<&J- ���ZAXS\UPR:LW�'CU�� k�$� | 
�/�/�/4�??j�&ELE�M/ T $1Uc c1j"NO�7�0�a3UTOOi�2H�A�4�� $DA{TA" T&e0   @P:�0� 2 
&PNP% ��P!U*.n   oFSyCjHrB� zB(�F�D(�1�R5C�DROBOT��H�CQBo�E�F�$CUR_"�B8�&SETU�	 �l� �P_MGN��INP_ASS � @�� �3�8"7�GP U�>VhSP!��&T1�
@B\8�8�T= 0 P�+ Kec1VRFY�8�T$5"&1� ��W��1�$R�/DSPH/ ([ �#A��#A�#A3tBOX/ 8�0������`bo%c4�TU�IR�0  ,�[ �62`ERa02� $k` ��a_S�bP�fZ}N/ 0 [9d&0� arZ_�  _� tu0  �@�A�Yv	�on ���$$CL,P  �����q��Q���Q�$' 2 ��uQ  G ��q���b0)�p�}�p��~ �4�F���m��� ���ǏُL����� ��E���i�{��� $�6��Z�����A� ��Ɵ؟��������2� �V�h�z�+���O�a� ԯ����
�@�Ϳ��� �v�'Ϛ����п^� �ϥ����<�N���r� �5�Gߺ�k����ϡ� �������\��ߒ� C��g�y��ߊ��"� 4���X�	����?��� ����������0��� T�f�x�)��M_�� ����>� t%���m\� ��:L�p� 3/E/�i/��q// �/�/�/Z/?~/�/A? �/e?w?�?�/�? ?2? �?V?OO�?*OOO�? �?�O�?�O�O.O�ORO dOvO'_�OK_]_�O�_ �O__�_<_�_�_r_ #o�_�_�_ko�_�o�o o�o8oJo�o�o1 C�og�o�o"� ��X	�|��� O�u�������0�� T���)���M���ҏ ��������,�ʟ�b� t�%���I�[�Ο�� ��ǯ:����p�!� ������i�ܯ�������$DCSS_C?SC 2I�ɱ�Q  D���@���&��� J�\�n�=ϒϤ϶υ� ��������"�4��X� j�|�Kߠ߲��ߓ��� �����0�B��f�x� ��Y���������� ���>�P�b�1������g�����������G�RP 2ɻ 	��	��cN� r����� �;&Kq\�� ����/�%// I/4/m/X/j/�/�/�/ �/�/�/?�/3??W? B?{?f?�?�?�?�?�? �?�?OOAO,OeOPO �O�O�O|O�O�O�O�O ___O_:_s_�_T_ f_�_�_�_�_o�_'o o7o]ooo>o�o~o�o �o�o�o�o�o5
�STAT 2�ɹY�,8���p�-�l��?b
?����XFL9C�/�?W�b?��=��D����D4��D����ɱ,p8xq?Y-��?����2t�4���?� � �q��p4��Z�C���CC����ɱxq��$����?]�˿�<h���������y�l��¤	~DcW���u�q��p9������ĸ�����|�˚��~� �=i�T�u��M@�=���?�~�^�p�,�Dq�?�,�X2N�=�N�DhBr�D�vD��E�X�ߺK=1�"�?~9���0�?X2K��N���W�e�����q��{��~́ɵ ��ɵ�J�\�:��� ���z�p�����uğ��؟�r��t��t ���bÒ�[Dc[���h�� t�������ԯ����� d��H�Z�8�~������䯺���ƿ��l����������M�' ����Z�� Vϐ�zόϮϰ�n�� ���>�P�.�t߆�d���p��s\�?a�܀���N�9D���X?���=�"�p�����D����|�*�p��t�x�l��t���p��{%��p���p��p6�����������n_4¤4�����92�ۤ��ǉ�p<���L��=�J�W�R�=���ih�Y�p�,�G��x�|�Z=�O_�DhA㈀���ꐇ�=1�~ꠀ�����W��kO�[����� ��߹���l�>�P�.� t���d������������������ ��(��0��4��b�>L��DcZ�2 ����� �� 0B��RxV�� ������� /������ۭ��׉��4��4�8��/./�/
/�/�/ �/�/�/",?>?�N? t?R?�?�?�?���� ���� ��$�6�H�Z� l�~���������O �?�? ��?l_~_\_�_ �_�_�_�_�
?o�/  oJo@RdvTo�o ho�o�o�o�o
�_ dvT����� �_6�J�B�,�J/ \/n/<�^�`���̏�� ���,�R\�n���� ����ȟڟ�?*_<_�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ��P_Ƛ��ҿ ��¿�� �:�D�� P�z�po�o�o�o���� `�����(�R�<��� �ߦ߄����ߺ� �� ,�f�<�B�H�r�h�z� ����|��������� �2�4��ߌ���|��� ������
��Z�l�*� <�N�`�r��������� ̯ޯ���&�8�J� 4F�������/ �/8/�H�j�l�F� �/�/�ϲ����ϴ/? �/"?L?6?X?�?t�J/ �?/�?�?�?�?0OBO \/�?lOr?xO�O��� ���O_�O_D_._ P_z_d_"O�_�_�_�_ o�_(o:ox��Z l~������ � 2DVhRo dovoo��o �2� �V�h�NO�_���_�� ȏ���/�/�/�F� 0�R�|�f������_� ��F��*��:�`�z� ��Ɵȟ����ү�O�O �O�Oܯ>���J�t�^� ����Пr��>���"�  ��X�jϨ���o �o�o�o�o��o ,>P�t��߂� �Ϧ�H��,�
�P�b� @���~������ ���� ��$���d�� `�����������x� $v�HZ8~��� ����������
� ��nXz�� �� 
//n@/R/ 0/b/�/f/���ߨϺ� ��������&�8�J� \�n߀ߒߤ߶��߲/ �/�ߘ/JO�/:O�O�O pO�O�O���O��O (_�0�B�T�2_�_F_ �_�_�_�_ o�_�OBo To2oxo�oho�o�o�O o�o�_�o 
(: L�>���� �
��o:�L��op����`�����Ƈ�$DC�SS_JPC 2��eQ G( D��Et� $�6�H��l�~���_� ��Ɵ�������ݟ2� D�V�%�z�����m�¯ ԯ毵�
�����R� d�3�������{�п� ��ÿ�*����`�r� AϖϨϺω������ ��&�8�J��n߀�O� a߶��ߗ�������� 4�F�X�'�|��]�o� �����������B� T�f�5�������}��� ������,��Pb tC������ ��(:	^p� Q����� // �6/H//)/~/�/_/ �/�/�/�/�/? ?�/@D?V?%?7?Cv؅S���@BS �HALT�?u5u? � Ip=����?�?�4�?�?O�6! O2ODO�6`OrO��O�6�A�O�O�O�3�O�OC_�6 _2_�_B�6`_r_�_�6	�_�P��_ox?Du�_Eo o*o{oNo�oro�o�o �o�o�o�o�oA& wJ\n���� ���=��a�4��� X�j�����ɏ���֏ �9���0���T�f� ����������ҟ�"� G��,�}�P���t�ů ������ί	��C�� (�y�L�^�p������� ��ʿܿ�?��$�b� ��Z�lϽϐ��ϴ�� ����;��I�2߃�V���?_MODEL ;2�;xt�i�W
 <m�c�:�H�J"����X�/�A� S�e�w������� ������+�=���a� s��������������� g�P��+�o� �������L #5�Yk}�� � /��6///1/ C/U/g/=�/a�/�/ ?�/�/D??-???�? c?u?�?�?�?�?�?�? �?@OO)OvOMO_O�O �O�O�O�O�O�O�/�/ �/__�_�Om__�_ �_�_o�_�_8oo!o 3oEoWoio�o�o�o�o �o�o�o�ojA S�;_M_{��u ����+�x�O�a� ����������͏ߏ,� ��b�9�K�]�o��� ������ɟ���� �p��Y�k������� �ůׯ$�����l� C�U���y���ؿ���� ӿ ���	�V�-�?ό� '�9�K�yϋ�a����� .���d�;�M�_�q� �ߕ��߹������� �%�7�I��m���� ������&������ ��E�W���{������� ��������X/A �ew���� ��B+=�� 7�ew���/� /P/'/9/K/�/o/�/ �/�/�/?�/�/�/L? #?5?�?Y?k?�?�?�? �?�O��?�?ZO1O CO�OgOyO�O�O�O�O _�O�OD__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o�?�o#OQo co�o�o�o�o�o %7�[m�� �����8��!� n�E�W�i�{�����uo ���oǏُF��/�|� S�e�w�ğ������џ �0���+�x�O�a� ������䯻�ͯ߯,� ������=�O��� 7�����ɿۿ�:�� #�p�G�Y�k�}Ϗϡ� ������$�����1� C�Uߢ�yߋ���s��� ����2���-�?�Q� c����������� ����d�;�M���q� ������������ N����);�#� ����&�\ 3EW�{��� �/��/X///A/ �/e/w/�/_q��/ �/�/??f?=?O?�? s?�?�?�?�?�?O�? OPO'O9OKO]OoO�O �O�O�O_�O�O�O�$��$DCSS_P�STAT ����cQQ?    t_�Z r_ (�_�_�WpkPkP�_�_ l cdP��P;_4oFo�)"ocUcUdovo�TTSETUP �	cYB�&T�#��!�dOYT1SC �2
�j`�!Cz��#/}�eCP [R�l�� DSo z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ��.h%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛ���������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� ����}����������� ����1CUg y������� 	-?Qcu��������Z�D �/*/</�/`/r/�/S/ �/�/�/�/�/??�/ 8?J??[?�?�?a?�? �?�?�?�?O"O�?FO XOjO9O�O�O/}O�O �OoO__0_�OT_f_ x_G_�_�_�_�_�_�_ �_o,o>ooboto�o Uo�o�o�o�o�o �o:L�O)�� ���� ��$�� H�Z�l�;�����q��� ؏ꏹ�� �2��V� h�z�I�������� ��_՟.�@�ǟd�v� ��W�����Я����� ��<�N��_����� e���̿޿����&� ��J�\�n�=ϒϤ�s���$DCSS_T�CPMAP  �������Q @ ~�J~�~�~���~�U~�~�~�	g�W  ~�~�~�U~�~�~�~�U~�~�~�~��~�~�~�~��~�~�~�~��~�~� ~�!~�"�~�#~�$~�%~�&�~�'~�(~�)~�*�~�+~�,~�-~�.�~�/~�0~�1~�2�~�3~�4~�5~�6�~�7~�8~�9~�:�~�;~�<~�=~�>�~�?~�@��UIR�O 2�����$��"�4�F�X� j�|��������������0�B�T�}� �}����������� ��1CUgy �����^���� �-?Qcu�� �����//)/ ;/M/_/��/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�?��?v/O��UIZNw 2��	 �����PObOtOy�KO�O �O�O�O�O�O_�O0_ B_T__x_�_�_k_�_ �_�_�_�_o,o�_Po boto�oIo�o�o�o�o �o�o:L^- ���i���� �$�6��Z�l�~�M� ����Ə؏�����ݏ�2�D�V�O��UFRwM R���� �џ���ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߒ��߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s��ߗ��� ��������'9 K]o����� ���#5GYk���x��� ���//�B/T/ //x/�/e/�/�/�/�/ �/�/?,??P?b?y ��?�?I?�?�?�?O O�?:OLO'OpO�O]O �O�O�O�O�O�O�O$_ 6__Z_l_�?�_�_A_ �_�_�_�_o�_2oDo ohozoUo�o�o�o�o �o�o�o.	Rd {_��9���� ���<�N�)�r��� _�������ޏ��ˏ� &��J�\�sw