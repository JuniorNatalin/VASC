A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �WVSCHD_T   H $FREQUENCY  $AMPLITUDE  $DWELL_RIGHT  $DWELL_LEFT  $L_ANGLE  �WVSCHDEXT_T  8 $ELEVATION  $AZIMUTH  $CENTER_RISE  $RADIUS  �8�$$CLASS  ������       �$WVSCH 2 ������� 
 ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  ?�  @�  =���=���B�  �$WVSCHEXT 2������� 
                                                                                                                                                                 �$WVSCHG  ������� 
                                         