��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�ASSNAME_�T   0 }$+ $'�WORD  ? L�EVEL  w$TI- OUTT� �&F/�� $SETUP�JPROGRAM�JINSTALL�JY  $C�URR_O�US�ER�NUM�S�TPS_LOG_ZP N��$�T��N�  6 CO�UNT_DOWN��$ENB_PCMPWD � �DV�IN!s$C� CRE�OPARM:� T:DIAG:)��LVCHK!F�ULLM0�YX=T�CNTD��MENU�AUT�O,�FG_DS�P�RLS����$$CL(   O���!��	���	�$DCS_C�OD@���%��  W'_S � *�! V&��A91("!�0 d $VA�G M/��R�J3ICSPEZ�VW���   5?67 TOR�$�#�P� ��!LINEBUILD�"?2007�%���� FANUC���25111�7 7��� B�EDIEN�%� 0O�&T �!J0�06�'  759�9���"6�&K=708;9608m;43J7D1�292�?10�:2]7�?011�%�� 9303�6�"�2�4^�38085�?1�7��14I5J4�923�5HG"G�154jO0�1:4�3653"O0�0�8003:4w1�G�4�D09�4J�FG� 118GF2��G�A36ZG(W�:5�97�O02J09q8�G(W6J425�_;02ZJ793�7(W�~J50Y(W�J416��G(W�J766�_0�2�J49}H(WZ4�93_032Z79%4o0�X�A1�_�`�J16_�`�[456B_03ZJ10�o�`�~J2�Y�g�J157�FO03�K29�o0�3�J734bo03vZ06�_J04�k�78�_04�;18v�o04J367��0�H�!�?�qZJ94�	h�w~J817�0l�h�Q85�04�J#13�8�w�K2)x�w�Z73�3�52Z54n�J10�:22UX ��J����6J����ZJ59H��N{䟊��J +����JO����Js��� Z�����5��Ǩ���`���֟��{50鏌_�ZJ43ŏ_�N{9��ȧ�J99��Ϡ�Lh��ȧ[7A_J11[c49�5-��:38���0��35J�1�[5�75Z�1�[����1�U���RyX0�r{�1i�0�λ86��1�QkL���1uk585~�1�k47E�`��;18�h`�J66���� ���qxX����^�J5c�C�q{9�iX��J3<o^�Rk8�_�Zq8[p���880�ߍ1%�82���J46��>�d�ZK������B���f�������
B�J4 �
��PDnp�ro�$�T��vE�G.!b#SU�!�n+�/�/b#WORD �!�9�n;�1
3�:d�,4 V�[t/&��jH �-4����