��   v��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<�$1_8k ���FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\9 ^75z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D��VCAX_�w A.  @ 5vFX0OR�@E ?NUM_SE238�_TO0Q�#RE_:� 2cT �+V>1 , $� �ME�vUPgDAT�wAXy_2 	8+VS5Q' 8<P��PnP;0k L\�R�PA�kQ�Q��+VM5Q  �$ISRTd 5+VG5Q { v��R2 
v�S2�T kR9�P 	��$U1SS  O����a����w�$' 1 �e� } �� 	 ����o�o�o�fт�p ������� `R�(a��o�oA,eP���xu}�a��|��:P[h#����9��.?4���|���n�|�+�=�d�a��V�s	� Q�w� 3Z� ��y�a�tB ��]��  ��B���f� ����������K��_������.���o�B������9�p�*pp���d�1�xC�U���=L��`�f��?�����@��� ͟ߟ���'�9�K�`]�o������� �eྯ̧��쯄d  2  ��/�A�S�e�w�����������<���� ��1�C�U�g�yϋ� �ϯ����`�a�o��� ���*�<�#�`�K߄� oߨߓ�c��ߡ���� &�[�5�G�n�k�}�� �����������"�� �P�b�t��������� ������(:�� ^p������E ϯ��6HZl ~�����˿� / /2/D/V/h/z/�/ �/�/�/�/���/��/ .??R?9?v?a?�?�? �?�?���?�?OO<O 'O�?]OoO�O�O�O�O 3O�O�O_�O_J_=� k_}_�_�_�_�_�_�_ �_oo1oCoUo|o �o�o�o�o�o�goio �o-#Tfx�� �������,� >�P�b�t��������� Ώ����/�(��L� 7�p�W������ʟ�� ��?�՟6�!�Z�l� �O{�������ïկQ� ���2�D�/�h�[_�� ������ѿ����� +�=�O�a�s�5�Ϭ� ��������G���'� K�Ar߄ߖߨߺ��� �������m�J�\� n�����������������$FMS_GRP 1^�� �>�IcsvGm��ZH�bI���+I��HH��O:J�Me%nO��<GN���J�^,3J��J����J�B�  ������4VA!��s�e3+�
��a�Ϝ�Cs��J���� N�he)P�L�O���xKP�K��K�{���o@��z?�z���Ict;Gm�#�H��[�_��H�P�+�Xk���(�����	p����3� �� 	W�7NQ;�W7O_W7P�G�G}�G�W7QWV:QWFW�W��W��Ui�<�V��V���W6^bX�,X�a���4�(�*�8���@�{C��A��;���A����o��EK��$!�q����e���Ra�6<� �!� ���� �� �K׏���M��X���|��-��J}�}����$�ƾ�������c�������4��R�_'M��������[�����7 �"^~ "G� �"2� "?� �"4h "� �"� !�k �!�� !һ �"�� # � �#� "����ܰ;�M �z zӖ zψ ��7��������>���҈������������<��������L����� <����w���1� �����a�9G� ���������a� R���(K�"4�W�4����4�q0:��4غ�4���4��4�)��4�
�4���1��1n��1��1?��:���dY��Ҳ������ҳ��2[o�7�ӧ��ӥ�[c0m�ӑ���ӓ��Ӗ?��ӗE�Ә��ә��Ӛ����t���o`���p���rC���8���:�����d����������}c"�}��3
�?�?�8�5R�4K|��3_��,�
�1��	��+�1��4��1_��_���4�"�	
�	��oED�)���[�_����
��26
4�{HwL��E�V�r_ж_��C[��WGu4�,����A�D�A
�_w���@_Ц_���_�V�A�*Q�_��
�T�%���T�A�WH2B@oI�	U�D.U4��P+_��_��_U�4��oo'o1f�5�1�p�4Yoko}o Wo*YFF�d+4�5�o�fE=4�;�h�a	�#�h�17���o������ф�����R���)������єʿ���8��y����n`�͏����ѿ͙п���c��6�����ܿN8�O� ?r�A�7?�#�?#�y?�#��?#�?�#��?#�Q?�#��?$�?�$w?$2�?�!�>?!�k?�!�!?"">�4�Z>�s>�ml>���p�k?V3�b�������5���� ��ձ�����p�6��E���#+��5ο��G<�������N���տ���W��E���I��2��w2{�r��T7��7���7����7��7����7���p��7����7�����7���:��#�T�:�w+�I���U�(������1�;��:�"��O���PsS� ���RB��N���Mۿ�H����E2��Cj���BJ��.����3�w���(����繿w5����Q��}#��O��^Or���?��?���?�߱?�ޣ?��z���᷀�?��p?���j?�|?�z�?�{"ˀ�@�v@#��?=]V?=Z}�X?��X	�,($MAKRO080�o'���4��UP022=�g�N� ��r��������̟	� ��?�&�c�J�\��� ������ɯ�گ��� ;�"�$�q�,�09���]�39�aÿ������ �π�)�S��w�b� �φϿϪ�������� �=�(�a�L߅ߗ�~� �ߦ������oY3� �oW�i�{����V��� R��������/�A�S� e�$���������~��� ����+=Oa  ����z�� �'9K]�� ��v����#/ 5/G/Y//}/�/�/�/ r/�/�/�/�/?1?C? U??y?�?�?,̫G�? �?�?�?i?"O4OFOXO O|O�O�O_O�O�O�O �O�O_0_B_T__x_ �_�_[_�_�_�_�_�f���1234567890o'e-�oIo 9omo]oyo�o�o�o�o �o�o�o!-5G {k������ ����S�C�_�g� y���������ӏ��� ��7�a���ﲟ ���ӟ���0�� T�?�x�c�u�����ү ������,�#�P��_ t�������	����o� ��(��L�^�pς� AϦϸ����ϛ� �� $���H�Z�l�~�=ߢ� �����ߗ���� ��� D�V�h�z�9����� �����
����@�R� d�v�5����������� ����<N`r 1����?�� 8J\n-� ������/� 4/F/X/j/)/�/�/�/ �/�/�/�/?oc�9? Q�]?M?i?q?�?�?�? �?�?�?OOO%O7O kO[OwOO�O�O�O�O �O�O�O_C_3_O_W_ i_�_�_�_�_�_�_�_ oo'oQoAouou�? �o�o�o�o�o�o  D/Aze��� ������@�7� d�v��/������Џ/� 􏃏�*�<�N��r� ����U���̟ޟ🯟 �&�8�J�	�n����� Q���ȯگ쯫��"� 4�F��j�|���M��� Ŀֿ迧���0�B� �f�xϊ�IϚ����� �ϣ���,�>���b� t߆�Eߖ߼������ ��(�:��^�p�� A�������� �� $�6���Z�l�~�=��� ���������� 2 )?MeoYas�� ����' [Kgo���� ����3/#/?/G/ Y/�/}/�/�/�/�/�/ �/�/?A?1?e?U?q?�y?�1�$PLCL�_GRP 1����1� �D�0�?��  �:[�?uض�9�O�:O%O ^OIO�OmOO�O�O�O �O _�O�>2_�OY_�O }_h_�_�_�_�_�_�_ �_o
oCo*o$_vo8o �o4o�o�o�o�o	 ?*cN�nho �|�x��)�� M�_�J���n�����ˏ�=�$VCAX_wREF�0 2�5� t 
 ����ERENCE 1��׏7�I�[�m�������2�ԟ���@
��.�@����3ß |�������į֯�S��4k�$�6�H�Z�l�~������5�̿޿ ���&�8ϣ���4 ��zόϞϰ���������7c��.�@�R�d�v߈����8����߀������0���9 ��l�~���������C�FACTOR?Y DATA\�� '�9�K�]�o������9������������	 ��GYk
�2_�����`����2_ �Pbt���� 'j�?�
//./@/ R/d/'���/�/�/ �/�/�/?'���/H? Z?l?~?�?�?�?'b� 7?�?OO&O8OJO\O '
��?�O�O�O�O�O �O_'�ՇO@_R_d_ v_�_�_�_'Z�/_�_ �_oo0oBoTo���_ �o�o�o�o�o�o�o�� /ASew% �����3�� %�7�I�[�m���_�t 7��Ώ�����(� �����d�v������� ��П;����/��0� B�T�f�x�㟥�/?�� Ưد���� ����� �?\�n���������ȿ 3���O��(�:�L� ^�p�ۿ��'_�Ͼ��� �����߃ϥ��_T� f�xߊߜ߮���_oqo ����,�>�P�b�t� �����������@�(�:�L����4� ��������������*� p���0BTfx� �S����  2D����� �����W�� (/:/L/^/p/�/�/� K��/�/�/??*? <?�/�x?�?�?�? �?�?�?O?�� O2O DOVOhOzO�O�?C� �O�O�O�O_"_4_�� ��j_|_�_�_�_�_�_ �_��	�o!o3oEoWo io��o�o�o�d