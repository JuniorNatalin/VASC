��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���F�SAC_LST_�T   8 �$CLNT_NA�ME !$I�P_ADDRES}SB $ACCN �_LVL  �$APPP   װ�$8 AO  O���z����w�$'DEF\ �w { �����ENABL�Ew �����L?IST 1 z�?  @!���������= "sF�j��� ��/�9///o/ B/�/f/�/�/�/�/�/ �/�/5???,?}?P? b?�?�?�?�?�?�?�? 1OOUO(OyOLO^O�O �O�O�O�O�O�O_ _ >_$_u_H_Z_l_�_�_ �W