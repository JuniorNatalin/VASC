��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���W�VSCHD_T �  H $F�REQUENCY�  $AMP�LITUDE@D�WELL_RIG�HTNLEF]L�_ANGLM&E�XT- 8 �$ELEVATI�ON@ZIMUT�H@CENTER�X SMRADIU�S@��$$C�LASS  �����������$' 2 ��� 
 �?�  @� =�{��B�  � "4FXj|�����  2� ���//+/=/O/a/���G  �� �/�/  