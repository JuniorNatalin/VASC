��  IL�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���S�BR_T   �| 	$SVMT�R_ID $R�OBOT9$GRP_NUM<AXISQ6K 6�NFF3 _PA�RAMF	$�  ,$MD �SPD_LIT�d&2*  �� � ���$$CLASS ? ������� � �$'  1 ���  T����R-200�0iB/185L���aiS�R30/3	 8�0A��
H1 DSP1-S1���	P01.03�,  	��  ��� � ��b���������
�=�#�r�9  ~��%����8 l��  ����x�� %��  ץ�� ����������  �2'-b��>���q�G�R����b���&��� �% ���� ͭ������������ �c6�����6N�������c�9	`B 0� �$  �� �:?p��@  'bx�'/�/�/�/L�/���/�/S�?)?;?  Z���2�'{�O��r�+� �3 ����=�����1�%m�>?L�?��� $J62@2HZ�l;���8�Ì��,p�@��n����o��o���#�q 3 ��|0����k)�2!�h	����u  �_��� u$t�?�4$��.>'���W
b����T'�`/r/�!d �/T_f_x_�_�/�_	?��_�_??Q? 3��2��<�����n	��0��4h� `z��1�`��D	��_Uo�?�?	�?63@BOKq m=R�3�IDONVL@��qI���keke�K^4�#����v�l���^7
���� �@�� U$V\o�E�_�>(��x��/	��MX=_*_ <_��)�;��__��_ p�����oˏݏ��x�no�o �`/12/4.43;e4@4�oZC ~b�q��a1|6O p�$0w�� (H������F�� ����_�����0�@���� Y$�'�4$���$>!V�A�q�/��������  ��������s~"��yO�ǯٯ���X�!��f(�M�_�q����������˿,�L�65@5p������ਗ�䴟ƟhArܑ
�a�� ��� �������+ ���>�Z$�������)�If���`���������������u� �ߙ߫����*���� �)�;�M�_�q��޿�� �66@6`(�:�L�Cc<C�l��~�ؕǺ���ϸρ�����F 
��>�\$'���� ���g�.���8��u/��f�@�R� d�-?Qc�߇�� �����)�;����A�<aPPgu		u�ao��� ��//,/>/P/b/ t/�/�/�/�/�/�/�/?<�?8?J?\?n? �?�?�?�?�?�?�?�3 n`
O���pO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_"?�_�_o o2o�DoVohozo�o�o�; � =�EXT�ENDED AXkIS-��q���4/5�� H� �� -ND��0.93'���  PG��r  H�X��������  �{�'�9~�5
���� Zp�l� �ܑt▂������� �,�c�	`� 7� (��t Z��	�! �_�q��������� ď֏�����0�B�T�*��(OO|�>O PObO�����*�<� N�`�r���������̯ ޯ���&�8��_\� n���������ȿڿ� ����?����Yϴ�Ɵ �Ϡϲ���������� �0�B�T�f�xߊߜ� ��������@���,� >�P�b�t����� ��*�<���`�rτ�L� ^�p������������� �� $6HZl ~��������  2DVhz�� ����0�B�
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?��?�?�?�?�? �?�?OO&O8O�� ��O���O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o h?0oBoTofoxo�o�o �o�o�o�o�oROdO �O�O�Ot���� �����(�:�L� ^�p���������ʏ&o � ��$�6�H�Z�l� ~������o0"̟F Xj2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v���䏬� ��п�����*�<� N�`ϼ�������� ������&�8�J�\� n߀ߒߤ߶������� ���"�4X�j�|� ������������� �zό�6������Ϝ� ����������, >Pbt���� ���N�(:L ^p�����&��  =�EX�TENDED A�XISh����aiS4/500�0 40Ak�H  DSP -~�P00.39�� 	�  o��Pm� H�X��q����ԯ  {n�C �9~�5
�� �p� ��l� l�_��tn�b� �/�/�/�/
??.?e��c	`�� 7 (�"t Z�� :?��j���!>?�?�?�?�?n��?�?OO'O9OKO0]OoO�O�O�X�J� �On�����_$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho �o�o�o�o�o�o�o 
.@,��O�O� �O�O������ *�<�N�`�r������� ��̏ޏ����po8� J�\�n���������ȟ ڟ���Zl��� �|�������į֯� ����0�B�T�f�x� ��������ҿ.���� �,�>�P�b�tφϘ� ����*i!/%/7/ I/[/m//�/�/�ߦ� �������� ��E?W? i?{?l�~����?�� ������� �2�D�V� h��O=�/���S�e��� ��	-?Qcu ������� );߿Mq�� �����//%/ ���=/�������/�/ �/�/�/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?UO/OAOSOeO wO�O�O�O�O�O-/_/ Q/�Ou/�/�/a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �oO�o�o�o#5 GYk}��O__ �3_E_��1�C�U� g�y���������ӏ� ��	��-�?�Q�c��o u�������ϟ��� �)�;�M���e�� ��˯ݯ���%� 7�I�[�m�������� ǿٿ����!�}�E� W�i�{ύϟϱ����� ����U���y�#ߝ��� ���ߛ߭߿������� ��+�=�O�a�s�� ��������;��� '�9�K�]�o������� ���E�7� [�m�5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �����/+�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO�mOO�O�O�O �O�O�O�O_!_}/�/ �/K_�/�/�/�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o cO+=Oas� �����;_m___ (��_�_]�o������� ��ɏۏ����#�5� G�Y�k�}������� ş�����1�C�U� g�y���������/� A�S��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�q�͟�� �Ϲ���������%� 7�Iߥ�ׯɯs���� ��������!�3�E� W�i�{�������� ������/���S�e� w��������������� cߕ߇�P�߽߅ ������ '9K]o��� ���7��/#/5/ G/Y/k/}/�/�/�/�/ !3�/Wi{C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O��O�O�O�O_ _)_;_M___q_�/�/ �/�_?'?9?oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E W�O{����� ����/��_�_�_ x��_�_����я��� ��+�=�O�a�s��� ������͟ߟ��_ �9�K�]�o������� ��ɯۯ�I�[��� ����k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������ ��	��-�?�Q�c�u� �ߙ���'����=�O� a�)�;�M�_�q��� �����������%� 7�I�[�m���ϣ��� ��������!3E W�����ߠ���� ��/ASe w������� //+/��=/a/s/�/ �/�/�/�/�/�/?? q�-?����?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�OE/__1_C_U_ g_y_�_�_�_�_?O? A?�_e?w?�?Qocouo �o�o�o�o�o�o�o );M_q�� �_�����%� 7�I�[�m���_o�_ ȏ#o5o���!�3�E� W�i�{�������ß՟ �����/�A�S�� e���������ѯ��� ��+�=�����U�Ϗ �󏻿Ϳ߿��� '�9�K�]�oρϓϥ� �����������m�5� G�Y�k�}ߏߡ߳��� ����E�w�i��� ��y���������� ��	��-�?�Q�c�u� ����������+��� );M_q�� ��5�'��K�]�% 7I[m��� ����/!/3/E/ W/i/{/���/�/�/�/ �/�/??/?A?S?e? ��}?�	�?�? OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_�/]_o_�_�_�_ �_�_�_�_�_om?�? �?;o�?�?�?�o�o�o �o�o�o1CU gy������ �S_�-�?�Q�c�u� ��������Ϗ+o]oOo �so�oM�_�q����� ����˟ݟ���%� 7�I�[�m������� ��ٯ����!�3�E� W�i�{��������� 1�C���/�A�S�e� wωϛϭϿ������� ��+�=�O�a߽��� �ߩ߻��������� '�9ǿ��c�ݿ� ����������#�5� G�Y�k�}��������� ������{�CU gy������ �S��w�@���u �������/ /)/;/M/_/q/�/�/ �/�/�/'�/??%? 7?I?[?m??�?�?�? #�?GYk3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�/�_�_�_�_�_ oo+o=oOoao�?�? �?�oOO)O�o '9K]o��� ������#�5� G��_k�}�������ŏ ׏�����{o�o�o h��o�o������ӟ� ��	��-�?�Q�c�u� ��������ϯ��O� �)�;�M�_�q����� ����˿ݿ9�K���o� ����[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱���� ������/�A�S�e� w����	ϳ�-�?� Q��+�=�O�a�s��� ������������ '9K]o�ߓ� �����#5 G����������� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??w-?Q?c?u? �?�?�?�?�?�?�?O asO����O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_5?�_o!o3oEo Woio{o�o�o�oO?O 1O�oUOgOyOASe w������� ��+�=�O�a�s��� ���_��͏ߏ��� '�9�K�]�o��o�o�o ��%����#�5� G�Y�k�}�������ů ׯ�����1�C��� U�y���������ӿ� ��	��-ω���EϿ� џ㟫Ͻ�������� �)�;�M�_�q߃ߕ� �߹��������]�%� 7�I�[�m����� ����5�g�Y��}Ϗ� ��i�{����������� ����/ASe w������� +=Oas� ���%���;�M�/ '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?�}?�?�?�? �?�?�?OO1OCOUO ��mO��/�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o�?Mo_oqo�o�o �o�o�o�o�o]O�O �O+�O�O�O��� �����!�3�E� W�i�{�������ÏՏ �Co��/�A�S�e� w���������M? �cu=�O�a�s��� ������ͯ߯��� '�9�K�]�o������ ��ɿۿ����#�5� G�Y�k�}�ٟ럕�� !�3�����1�C�U� g�yߋߝ߯������� ��	��-�?�Qﭿu� ������������ �)��Ϸϩ�S����� �Ϲ�������% 7I[m��� ����k�3E Wi{����� �C�u�g�0/����e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?OO 'O9OKO]OoO�O�O�O //�O7/I/[/#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�?�o�o�o�o�o �o	-?Q�O�O �O{�O__��� �)�;�M�_�q����� ����ˏݏ���%� 7��o[�m�������� ǟٟ����k�� X���������ïկ �����/�A�S�e� w���������ѿ�?� ���+�=�O�a�sυ� �ϩϻ���)�;���_� q���K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������� ��������1�C�U� g�y�����ϣ��/� A�	-?Qcu ������� );M_��� �����//%/ 7/�������/�����/ �/�/�/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OgOAOSOeO wO�O�O�O�O�O�O�O Q/c/_�/�/�/s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o%O�o�o#5 GYk}���O/_ !_�E_W_i_1�C�U� g�y���������ӏ� ��	��-�?�Q�c�u� ���o����ϟ��� �)�;�M�_���� ����ݯ���%� 7�I�[�m�������� ǿٿ����!�3Ϗ� E�i�{ύϟϱ����� ������y���5߯� ��ӯ�߭߿������� ��+�=�O�a�s�� ����������M�� '�9�K�]�o������� ����%�W�I���m�� ��Yk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/���/+=? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[O�mO�O�O�O �O�O�O�O_!_3_E_��$�$SBR2 �1�%qP T?0 � �/�) �_�_�_�_�_�_o o,o>oPoboto�o�o {_�_�o�o�o( :L^p���� �o�o�o ��$�6�H� Z�l�~�������Ə؏ ����2�D�V�h� z�������ԟ��� 
����@�#�d�v��� ������Я����� *�<�N�1�r�U����� ��̿޿���&�8� J�\�nπ�c�L_���� ��������,�>�P� b�t߆ߘߪ߸ٚ��� �����"�4�F�X�j�|��������� ����#�5�G� Y�k�}����������� ������0BTf x������� ,>��bt� ������// (/:/L/^/p/T�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�/�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O�? �O
__._@_R_d_v_ �_�_�_�_�_�_�_o �O*o<oNo`oro�o�o �o�o�o�o�o& 
oo\n���� �����"�4�F� X�<h�������ď֏ �����0�B�T�f� x���n�����ҟ��� ��,�>�P�b�t��� ������������ )�;�M�_�q������� ��˿ݿ�"�$�6� H�Z�l�~ϐϢϴ��� ������� ߤ�D�V� h�zߌߞ߰������� ��
��.�@�R�6�v� ������������ �*�<�N�`�r���د ����������' 9K]o���� j����"4F Xj|����� ���//0/B/T/f/ x/�/�/�/�/�/�/�/ ?�?>?P?b?t?�? �?�?�?�?�?�?OO (O:O?^OpO�O�O�O �O�O�O�O __$_6_ H_Z_l_PO�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�_�o�o�o �o
.@Rdv ������o�� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�� X�j�|�������į֯ �����0�B�T�f� J���������ҿ��� ��,�>�P�b�tφ� j�|����������� (�:�L�^�p߂ߔߦ� �ߜ����� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
 �@Rdv ������� *<N2r�� �����//&/ 8/J/\/n/�/d�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�/�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�? __,_>_P_b_t_�_ �_�_�_�_�_�_oo �O:oLo^opo�o�o�o �o�o�o�o $6 o,ol~���� ���� �2�D�V� h�Lx�����ԏ� ��
��.�@�R�d�v� ����~���П���� �*�<�N�`�r����� ����̯�����&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0��T�f� xߊߜ߮��������� ��,�>�P�b�F߆� ������������ (�:�L�^�p�����x� �������� $6 HZl~���� ���� 2DV hz������ ��/./@/R/d/v/ �/�/�/�/�/�/�/? ?�(?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO.?nO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_`O�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�_�o�o�o ,>Pbt� ������o�� (�:�L�^�p������� ��ʏ܏� ���6� H�Z�l�~�������Ɵ ؟���� �2�D�(� h�z�������¯ԯ� ��
��.�@�R�d�v� Z�������п���� �*�<�N�`�rτϖ� z�����������&� 8�J�\�n߀ߒߤ߶� �߬������"�4�F� X�j�|�������� �������0�B�T�f� x��������������� ,�Pbt� ������ (:L^B��� ���� //$/6/ H/Z/l/~/�/t�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�/�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O�? _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 
_Jo\ono�o�o�o�o �o�o�o�o"4F *o<o|����� ����0�B�T�f� x�\������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ�� ��$�6� H�Z�l�~�������ƿ ؿ�����2�D�V� h�zόϞϰ������� ��
��.�@�$�d�v� �ߚ߬߾�������� �*�<�N�`�r�Vߖ� �����������&� 8�J�\�n��������� ��������"4F Xj|����� ���0BTf x������� ��,/>/P/b/t/�/ �/�/�/�/�/�/?? (?/8?^?p?�?�?�? �?�?�?�? OO$O6O HOZO>?~O�O�O�O�O �O�O�O_ _2_D_V_ h_z_�_pO�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�_�o�o *<N`r�� ������o�&� 8�J�\�n��������� ȏڏ����"�4�