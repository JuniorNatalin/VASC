A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DCSS_CPC_T   � $COMMENT $ENABLE  $MODE  $GRP_NUM  $MODEL_NUM   $UFRM_NUM  $NUM_VTX  $X   $Y   $Z1  $Z2  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD  �DCSS_CSC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $TCP  $UFRM_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  �DCSS_GRP_T  � $TCPCHG_SIZE  $APSPD_MODE  $ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $APSPD_JMODE   	$ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$TCP_SEL  � �DCSS_GSTAT_T  D $FP_BASE $LINK_BASE ! 	$LINK_BASE_V ! 	$LINK_BASE_H ! 	 (�DCSS_JPC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $UPR_LIM  $LWR_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD   ��DCSS_JSC_T  | 
$COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  ��DCSS_ELEM_T  T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    "D�DCSS_MODEL_T   $COMMENT $ELEM 2 
�DCSS_PSTAT_T  � 	$STATUS_CPC    $STATUS_CSC   $STATUS_JPC   ($STATUS_JSC   ($USER_MODEL   $ROBOT_MODEL   $USER_ELEM   $ROBOT_ELEM   $CUR_TCP   t�DCSS_SETUP_T 	 l $DISP_MGN  $INP_ASSIST  $TOOLCHG_ENB  $DO_TYP  $DO_IDX  $DO_MGN  $CALMD_ENB  $CALMD_STAT  �DCSS_T1SC_T 
  $ENABLE  $SPD_LIM  �DCSS_TCP_T  l $COMMENT $UTOOL_NUM  $MODEL_NUM  $VRFYIO_TYP  $VRFYIO_IDX  $X  $Y  $Z  $W  $P  $R  X�DCSS_SPH_T  ( $SIZE  $DATA1  $DATA2  $DATA3  �DCSS_BOX_T  8 $SIZE1  $SIZE2  $SIZE3  $X  $Y  $Z  $R  ��DCSS_TUIRO_T  , $TYPE  $SPHERE 2 $BOX $BOX_S 2 ��DCSS_TUIZN_T  0 $ENABLE  $X   $Y   $Z_UPR  $Z_LWR  �DCSS_UFRM_T  @ $COMMENT $UFRM_NUM  $X  $Y  $Z  $W  $P  $R  t�$$CLASS  ������   Q    Q�$DCSS_CPC 2 ������Q   ��                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �$DCSS_CSC 2������Q  D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_GRP 2������Q  �                         	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                         �$DCSS_GSTAT 2������Q  ,8��p�:>��0�N�>��?q����=�(��rh�|:oD���D�<KDBy���� 	 88�?D`?$��    �X�|4�j?�  ?$�ݿD`4��ZCo]CH��    ���8�>�&;>a!�?p�n�8G���0>��?$�ݿD`4��ZD*�C�rlD|�����8�><=�|?|�$��?D]��CL�A o�"�>1מD	�uC��D������8�<��N>x�I?xG��A r�"�>1ך?'��<*K>/'D���D��D|\\���8�?? ?*db�+�%�'��?<*L�/��(�>rS?|:oD���D��D|\\���8��p�:>��0�N�>��?q����=�(��rh�|:oD���D�<KDBy����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX��� 	 88�?Di?$��    �X�n4�p?�  ?$�ҿDi4��ZCohCH��    ���8�>�&+>a!Q?p�s�8G���)>��?$�ҿDi4��ZD*�C�rHD|�����8�>;/=��?|�$��?Df��C}�A ��"�>1�vD	�bC�QD������8�<��>xɤ?xG��A ��"�>1�r?'�տ<*[>/OD���D��D|\����8�??)?*dW�+y>�'��?<*\�/:��*x>q�?|:mD���D��D|\����8��p�,>��W�OH>��8?q������=�*j�qܿ|:mD���D�<?DBzX���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8�����������������������������������������$DCSS_JPC 2������Q ( D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_JSC 2������Q ( @BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                               =���BS HALT                                               =���BS HALT                                 	              =����                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �$DCSS_MODEL 2������Q x�                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �$DCSS_PSTAT ������Q       (  (     ����                                                                                    ������������                  �������������$DCSS_SETUP 	������QB�                B�          �$DCSS_T1SC 2
������Q      Cz      Cz      Cz      Cz      Cz      Cz      Cz      Cz  �$DCSS_TCP R������Q � 
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �$DCSS_TCPMAP  ������Q @                            	   
                                                                      !   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @�$DCSS_TUIRO 2������Q �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$DCSS_TUIZN 2������Q 	 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �$DCSS_UFRM R������Q � 	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      