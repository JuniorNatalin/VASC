A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DMR_GRP_T  � $MASTER_DONE  $OT_MINUS   	$OT_PLUS   	$MASTER_COUN   	$REF_DONE  $REF_POS   	$REF_COUNT   	$BCKLSH_SIGN   	$EACHMST_DON   	$SPC_COUNT   	$SPC_MOVE   	$ADAPT_INER   	$ADAPT_FRIC   	$ADAPT_COL_P   	$ADAPT_COL_M   	$ADAPT_GRAV   	$SPC_ST_HIST   	$DSP_ST_HIST   	$SHIFT_ERROR  $SPC_CNT_HIS   	$MCH_PLS_HIS   	$ARM_PARAM   d$MASTER_ANG  $DSP_ST_HIS2   	$CLDET_CNT   	$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$GRAV_MAST   ,�FMS_GRP_T t *$REM_LIFE   	$NT_LIFE   	$T_LIFE   	$CLDET_ANG   	$CLDET_DSTB   	$NT_LIFE_0   	$T_LIFE_TEMP   	$REM_LIFE_0   	$GRP_CL_TIME  $PCCOMER_CNT   	$FB_COMP_CNT   	$CMAL_DETECT   	$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $DTY_STR_T  $DTY_END_T  $CLDET_CNT   	$CLACT1   $CLACT2   $CLACT3   $CLACT4   $CLACT5   $CLACT6   $CL_OVR   $CLOMEGA1   $CLOMEGA2   $CLOMEGA3   $CLOMEGA4   $CLOMEGA5   $CLOMEGA6   $CL_FRMZ   $CLDEPT_IDX   $CLCURLINE   $CLDEST1   $CLDEST2   $CLDEST3   $CLDEST4   $CLDEST5   $CLDEST6   $CLNAME ?( �PLCL_GRP_T  � 	$CALIB_STAT  $TRQ_MGN   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	��VCAX_REFA_T  @ $REF_FACTORY  $NUM_SET  $MAST_TO_REF  $PRE_MST2REF   ��VCAX_REFD_T  , $COMMENT $REF_UPDATE  $REF_AXIS 2 	��VCAX_REFS_T  8 $STEP_MS_ENB  $NUM_SET  $STEP_DATA  $PRE_STEP  �VCAX_REFM_T   $IS_SET  $MASTER_COUN  �VCAX_REFG_T  0 $REF_DATA 2 
$REF_STEP 2 	$PRE_MASTER 2 	�$$CLASS  ������       �$DMR_GRP 1 ������      	                                      	                                      	  �� :���Y4�   �O s�;                	                                      	                                      	                                 	                                	  1:� �09�)����������             	                                      	                    	                    	                    	                    	 ��������2��       	    ��         	 B  B B   B  B                  	  i4EKt ��6I�v�R j�             	 �?�0��� �3��D �2� u#�             d                                                                                 =L��                                    ?�                              @�                                                                                                                                                                                                                                                           	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                         	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 ����    	                                      	                                      	                                          	                                      	                                      	                                      	                                     	                                      	                                      	                    	                    	                    	                    	                    	                    	                                          	                                      	                                      d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                             	 ��������������������������� 	 ���������������������������     2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                 �����$FMS_GRP 1������  	 KkF�H��H
��K��J��	I���             	 LKZOS�O�<�I�$:J`<yI��6             	 B�  B�  B�  B�  B�  B�               	 AgjH�_��A�[w
¢DDB���             	                                      	 M���P���Q�JK!�9K���J��             	 AбiAбiAбiAбiAбiAбi             	 KkF�H��1H
��K��J��I��7            W7� 	                                     	                                      	                                                                              Vϱ�V�7V�DVӈ�VԭV՘�V՚�V՜Vա�W7cW7uW7zW7�W7�W7�VȀRVɄ�VɅ V̲OV�<Xӭ�Xհ� 	       
             +              ���J��̊���u���s��˧�����������m���} C�u C�[ C�G E1� E�� Fn����N�������K�����ː  �u\$�uJG�uK�u\v�uP��u_%�uN��uPp�uO�-�g-/9-;�"�!�!��uHi�u`t�uN��uL��u3~   �5J �q� �nm �6� �h? �0M �gM �g� �j��z���y�|�z~�e���e$��d5� �v] �/ �g� �kj ���  �r��r��r�$�r�<�r�/�r��r��r���r� ]B� ]f{ ]Dz \� ^�) a�]�r���r��r���r�Q�r�(  ������\������C���x�����{S���v��#����������H�D  (�D(σ(��(��(ϲ(�/(�J(��(��%��%��%���dY���(Ѐ(�,(�(З(��     d   d   d   d   d   d   d   d   d   
   
   
   
   
   
   d   d   d   d   d  ���j�����������`�������������������    ����   ����   �������A���������������    P   g   �  Q   ,  �   K   L   '   ����               �  w   S      �  �����������������Y������������������G   ����      ���O���)������A����  ������V����������C���:��� ���B�����������   ����    �����������������������  �����������8�������������������l����                    ���p�������U������/  ���=���"���������1���A��� ��� ���   ��������          �������������������     d   d   d   d   d   d   d   d   d  -  -  -  -  -  -   d   d   d   d   d                                                            �                         "   "   "   "   "   "   "   "   "                     "   "   "   "   "  �3b�0G�0G�3b�0G�3b�0G�0G�0G>x�9>x��>u�P>}��>T|>�?�0G�3b�0G�0G�0G  >�}>��p>��o>�}>��p>�}>��m>��m>��p������ҿ��z1�z�Ŀy�[>��p>�z>��m>��o>��p  ��׾˛F�˛F��׾˛F��׾˛D�˛D�˛F>�Ɍ>�0 >�Bc>ߖP>��>��پ˛F��־˛D�˛F�˛F  �I���I�y�I�y�I���I�y�I���I�x�I�x�I�y���K���˿��� _��4��b��I�y�I���I�x�I�y�I�y  ?��?�Y?�Y?��?�Y?��?�Y?�Y?�Y��h#���M��h���z=���M��@�?�Y?��?�Y?�Y?�Y  @=.�@=,�@=,�@=.�@=,�@=.�@=,�@=,�@=,�?���?�\�?��3?���?��|?���@=,�@=.�@=,�@=,�@=,�  ,($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP006                                     ($UP006                                     ($UP006                                     ($UP006                                     ($UP006                                     ($UP006                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                     ($UP007                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456       	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                          	                                      	                                      	                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ,($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      ($123456789012345678901234567890123456      �$PLCL_GRP 1������� D    	 ?�  ?�  ?�  ?�  ?l��?qP"?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                          	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$VCAX_REF_GR 2������ t 
 �REFERENCE 1        	                                                                                                                                                 REFERENCE 2        	                                                                                                                                                 REFERENCE 3        	                                                                                                                                                 REFERENCE 4        	                                                                                                                                                 REFERENCE 5        	                                                                                                                                                 REFERENCE 6        	                                                                                                                                                 REFERENCE 7        	                                                                                                                                                 REFERENCE 8        	                                                                                                                                                 REFERENCE 9        	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE2_1       	                                                                                                                                                 REFERENCE2_2       	                                                                                                                                                 REFERENCE2_3       	                                                                                                                                                 REFERENCE2_4       	                                                                                                                                                 REFERENCE2_5       	                                                                                                                                                 REFERENCE2_6       	                                                                                                                                                 REFERENCE2_7       	                                                                                                                                                 REFERENCE2_8       	                                                                                                                                                 REFERENCE2_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE3_1       	                                                                                                                                                 REFERENCE3_2       	                                                                                                                                                 REFERENCE3_3       	                                                                                                                                                 REFERENCE3_4       	                                                                                                                                                 REFERENCE3_5       	                                                                                                                                                 REFERENCE3_6       	                                                                                                                                                 REFERENCE3_7       	                                                                                                                                                 REFERENCE3_8       	                                                                                                                                                 REFERENCE3_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                          
 �REFERENCE4_1       	                                                                                                                                                 REFERENCE4_2       	                                                                                                                                                 REFERENCE4_3       	                                                                                                                                                 REFERENCE4_4       	                                                                                                                                                 REFERENCE4_5       	                                                                                                                                                 REFERENCE4_6       	                                                                                                                                                 REFERENCE4_7       	                                                                                                                                                 REFERENCE4_8       	                                                                                                                                                 REFERENCE4_9       	                                                                                                                                                 FACTORY DATA       	                                                                                                                                                  	                                                                                                                                         	                                                                         