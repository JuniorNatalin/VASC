��   ?�A��*SYST�EM*��V8.2�306 4/2�
 014 A �
  ���M�N_MCR_TA�BLE   �� $MACRO�_NAME �%$PROG@E�PT_INDEX�  $OPE�N_IDaASSIGN_TYPD � qk$MO�N_NO}PRE�V_SUBy a �$USER_WO�RK���_L� M�S�*RTN � D&SOP_�T  � �$�EMGO���RESET�MsOT|�HOLl���12�ST{AR PDI8GU9GAGBGC��TPDS�RELt�&U� �� �EST���/SFSP�C��`�C�C�NB�B�S)*$8*$3%)T ''5%)6%)7%)|S�PNSTRz�"D�  �$$C�Lr   ��i��!�����:�LDUIMT  ��������$MAXDRI�� ���%
�$.1� �% �� d%Ope�n hand 1�����%ZG_M�ENUEC?��^�x3�!�?�a  %Close3?�F=�?�?���"  ��!�#S0CUST_MN �?I:�6&O�q:�6�l�w �8d 23O�OoO8O�3���UB�9eO�?�O�?�3��1�3Relax��O�OK_]_�9�6 __�_H_�_�=�"�1`�_�_�_o�_ �_ VoI:No�o�7�3Fo�o jo�o�o�o�o'�oK �o�0�Tf� �����G��W� }�,�>���b�׏���� ���
�C���y�(� ��L�^����П	��� ʟ?��c��$�^��� Z�ϯ~������)�د �$�q� ���D�V�˿ z�ۿϰ�¿7��[� 
�ϑ�@ώ���vψ� �Ϭ�!�����/�i�T� ��<�N���r��ߖߨ� ��/���S����8� ��\�n�������� ��O���_���4�F��� j���������K ���0�Tf� ����G�k ,f�b��� /�1/��,/y/(/ �/L/^/�/�/�/	?�/ �/??�/c??$?�?H? �?�?~?�?O�?)O�? �?7OqO\O�ODOVO�O zO�O�O�O�O7_�O[_ 
__�_@_�_d_v_�_ �_�_!o�_�_Woogo �o<oNo�oro�o�o�o �oS�8 �\n����� �O��s�"�4�n��� j�ߏ�����ď9�� ��4���0���T�f�۟ ������ҟG���k� �,���P���ׯ���� ���1���?�y�d� ��L�^�ӿ�������� �?��c��$ϙ�H� ��l�~ϸ�ߴ�)��� ��_��oߕ�D�V��� z��ߞ߰�%���"�[� 
���@��d�v��� ����!�����W��{� *�<�v���r������� ��A��<�8 �\n���� �O�s"4�X ����/�9/� �G/�/l/�/T/f/�/ �/�/�/�/�/G?�/k? ?,?�?P?�?t?�?�? O�?1O�?�?gOOwO �OLO^O�O�O�O�O�O -_�O*_c__$_�_H_ �_l_~_�_o�_)o�_ �__oo�o2oDo~o�o zo�o�o�o%�oI�o 
D�@�dv� ��!���W��{� *�<���`���珖��� �̏A����O���t� ��\�n�㟒����ȟ �O���s�"�4���X� ͯ|���ȯ�į9�� ��o�����T�f�ۿ ��������5��2�k� �,ϡ�P���tφ�������1�����
Se�nd Event�7��SENDEgVNTs��(K�� %	_�Datya��z�DATA��ڡ�'��%_�Sy�sVar��|�SY�SV;��)�%�Get��<�GE�T��d�*w�%R�equest M�enu���REQOMENU���+�� !�b�߆�A��ϼ�k� ��������(��L�� �1�gy� ���HZE~ -?�c����  //D/�/z/)/�/ M/_/�/�/�/
?�/�/ @?�/d?v?%?_?�?[? �??�?O�?O<O�? �?rO!O�OEOWO�O�O �O_�O�O8_�O\__ _W_�_�_�_w_�_�_ �_"o�_�_ojoo�o =oOo�oso�o�o�o�o 0�oT�9� �o������ P�b�M���5�G���k� ������ۏ(��L��� ���1���U�g���� �����ӟH���l�~� -�g���c�د����� ���D���z�)��� M�_�Կ�ѿ
Ϲ�˿ @��d��%�_Ϭϗ� ��ϑ�ߵ�*������%�r�!ߖ�E�W��$�MACRO_MA�X�������Ж��SOP�ENBL �������y�T�T��#����PDIMS�K���� �;�S�UE�W�TPDSB�EX  �S�U���߿�P�����