A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �PMC_CFG_T   � $PMC_NUM_MSK  $EXE_TYPE  $MEM_OPT  $MN_CNF  $IF_CYC_NUM  $IF_SCN_TIME  $RESET_PTIME  $CYCLE_TIME  $CHECK_DSBL  $DRAM_MARGIN  $STORE_TYPE     �PMC_DEV_T  d 	$PMC_NO  $PMC_CHAR  $PMC_ADDR  $SIZE  $RACK  $SLOT  $MOD_TYPE  $IO_TYPE  $OCCPY  �PMC_IF_T  L $PMC_NO  $PMC_CHAR  $PMC_ADDR  $PMC_SIZE  $IO_TYPE  $IO_IDX   ��PMC_TYPE_T  � 
$PMC_SEQ  $MEM_TYPE  $EXE_RATE  $CTR_TYPE  $BUFF_SIZE  $PMC_SIZE  $RUN_STATUS  $CUR_TIME  $MAX_TIME  $MIN_TIME    ��SNP_PARAM � $CHANNEL  $CONNECTION_  $CPU_ID   $BAUD_RATE  $NOISY_CHANN  $T1  $T2  $T3  $T3_PRIME  $T4  $MAX_DATA_SI  $QUEUE_DEPTH  $COMM_BUF_SI  $MAX_RETRIES  $AUTO_START  $PMC_TYPE  $BG_STORE  $DISP_INFO  $CYCLE_PMC  $LIMIT_PMC  $LAD_EXEC  $EXE_CYCLE1  $EXE_CYCLE2  $EXE_CYCLE3  $EXE_CYCLE4  $LAD_PRI1  $LAD_PRI2  $LAD_PRI3  $LAD_PRI4   |�$$CLASS  ������       �$PMC_CFG  �������                      d               �$PMC_DEV 2������� d $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$PMC_IF 2������� P       X       �            X  �      !         X  �               X  �               X  �               X                  X        !   )      Y       �            Y  �      "         Y  �               Y  �               Y  �      	         Y                  Y        "   )      F       �            F   �   �            F  �               F  �   ����         G       �            G   �   �            G  �               G  �   ����         K            '      K  �        '�      R      �     *�      D      �     '      G      H      A      F      H      A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$PMC_TYPE 2�������  (        d        �|                                                                                                                                                                                                       �$SNP_PARAM �������                                   �  '  '                                   U   d                            