A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �PASSNAME_T   0 $NAME $PASSWORD  $LEVEL  $TIME_OUT  ��PASSWORD_T � $SETUP  $PROGRAM  $INSTALL  $TIME_OUT   $CURR_LEVEL   $CURR_USER   $NUM_USERS  $PS_LOG_EVEN   $LOG_EVENTS  $LEVELS   $COUNT_DOWN   $ENB_PCMPWD  $DVPCM_LOGIN  $CALL_PCMCRE   $PARM_PCMCRE   $STAT_PCMCRE   $DIAG_PCMCRE   $PCM_LOGIN   $ENB_LVCHK  $ENB_FULLMN  $ENB_TIMEXT  $ENB_CNTDWN  $ENB_MENU  $AUTOLOGIN  $ENB_CFG_DSP  $ENB_RLS_DSP  8�$$CLASS  ������   	    	�$DCS_CODE  �   ���   	�  W�$DCS_CODE_S  ������   	�  �������������$PASSNAME 1 ������	� d $VAG MIN       RJ3ICSPEZVW        567 TOR        567 PER      ��  LINEBUILDER   2007LINEBUIL     FANUC         251117 7         BEDIENER      2010OPER           J006           7599               56 7           567                J008           6087               J009           7292               J010           6272               J011      ���  9303      �����    J012      ���  8085      �����    J013      ���  9499      �����    J014      ���  2313      �����    J015      ���  9543      �����    J016      ���  6535      �����    J017      ���  0036      w���    J018      ���  6090      �����    J019      ���  1182      �����    J020      ���  0364      �����    J021      ���  5973      �����    J022      ���  0988      �����    J023      ���  4258      �����    J024      ���  7931      �����    J025      ���  5020      �����    J026      ���  4166      �����    J027      ���  7668      �����    J028      ���  4915      �����    J029      ���  4932      �����    J030      ���  7946      �����    J031      ���  0188      �����    J032      ���  1682      �����    J033      ���  4454      �����    J034      ���  1082      �����    J035      ���  2023      �����    J036      ���  1579      �����    J037      ���  0298      �����    J038      ���  7345      �����    J039      ���  0620      �����    J040      ���  7781      �����    J041      ���  9186      �����    J042      ���  3675      �����    J043      ���  5303      �����    J044      ���  9426      �����    J045      ���  8171      �����    J046      ���  4859      �����    J047      ���  1311      �����    J048      ���  6234      �����    J049      ���  7918      �����    J050      ���  5420      �����    J101      ���  2221      �����    J102      ���  2221      �����    J103      ���  2221      �����    J104      ���  5912      �����    J105      ���  2221      �����    J106      ���  2221      �����    J107      ���  2221      �����    J108      ���  2221      �����    J109      ���  2221      �����    J110      ���  2221      �����    J111      ���  2221      �����    J112      ���  2221      �����    J113      ���  2221      �����    J133      ���  5059      �����    J134      ���  4371      �����    J135      ���  2909      �����    J117      ���  9971      �����    J118      ���  6044      �����    J119      ���  1764      �����    J120      ���  4972      �����    J121      ���  3804      �����    J122      ���  2352      �����    J123      ���  5755      �����    J124      ���  1239      �����    J125      ���  1122      �����    J126      ���  1150      �����    J127      ���  9865      �����    J128      ���  2219      �����    J129      ���  5853      �����    J130      ���  4749      �����    J051      ���  9830      �����    J052      ���  6601      �����    J153      ���  7736      �����    J131      ���  2345      �����    J132      ���  5555      �����    J136      ���  9031      �����    J137      ���  3668      �����    J138      ���  4881      �����    J139      ���  8202      �����    J140      ���  8800      �����    J141      ���  8249      �����    J142      ���  4636      �����    J143      ���  2221      �����    J144      ���  2221      �����    J145      ���  2221      �����    J146      ���  2221      �����    J147      ���  2221      �����    J148      ��  2221       ����    J149         2221      ��P��    npro       �  3579      EG.��  �$PASSSUPER  ������	�VAG MIN       RJ3ICSPEZVW      �$PASSWORD ������	��              �              �                                                                     d       V�[t&��j                                                                                                    