��  	��A��*SYST�EM*��V8.2�306 4/2�
 014 A�5  ����A�AVM_WRK_�T  � �$EXPOSUR�E  $CAMCLBDAT@ �$PS_TR�GVT��$X� aHZgDIUSfWgPgRg�LENS_CEN�T_X�YgyO�Rf   $C�MP_GC_�U�TNUMAPRE_MAST_C�� 	�GRV_}M{$NEW���	STAT_R�UNARES_E=R�VTCP6� %aTC32:dXSM�&&�#�END!ORGBK!SM��3!�UPD��ABS�; � P/   $PARA� �  ���ALRM_REC�OV�  � A�LM"ENB���&ON&! MDG�/ 0 $DEBUG1AI"d�R$3AO� TYPsE �9!_IF�� D $ENwABL@$L�T P d�#U�%Kx!;MA�$LI"��
 �APC�OUPLED�� $!PP_PR�OCES0s!�(1�s!"PC> Q�� � $SOF�T�T_ID�"TOTAL_EQs 3$0'0NO*2U �SPI_INDE�]?5X�"SCRE�EN_NAMr ��"SIGNe0��/�+!0PK_FI�� 	$THK�Y�7PANE24 �� DUMMY1�d�4d!�54�1_P�ARG�R�� � $TI=T�!$I��N �DdDd D�0D5��66�67�68�69�70�7G�1EG�1TE0G1:G1DG1NG�1XG2cB��A�SBN_CF>"� 8F CNV_J� ; �"L A_CM�NT�$FLA�GS]�CHEC��8 � ELLSE�TUP 	 P�� HOME_IO�z0� %5SMAC{ROARREPRJX{0D+>0�dR{lT���AUTOBA�CKU�
 }�)DEVIC�3TIc0�� 0�#���PBS$INT�ERVALO#IS�P_UNI��P_�DO�V7�YFR_F\0AINz1��x1�S�C_WA�T��Q-jOFF_� N��DELZhLOGp�R�1ea�R?�Q�f`�3?�� {1�5�ϴ�MO� ZcE D [MZc����aREV�BIL~�gt�AXI� ~�bR  � �OD7P�a$�NO�@M���cr�"w� �u<q XZ0D~�C d E �RD_E�`Ts �$FSSBn&$CHKBD_SE�U�AG G�0 ?$SLOT_�V2�q� Vzd�%����Q_EDIm  � � cQG��CPS:`a4%$�EP1T1$OP�^02dap_OKvnrUS�!P_C� ��q�T�vU UPLACI4!TQ?��p( �Q�COMM� e0$D;�Q�J0f`�y�?�2���BL%0OU�r ,K�QQ2QU B�@y O]Å���CFWt X $GR� ��{MBZ`NFLI�<��0UIRE��$�g"� SWITCH^��AX_N)PSs"�CF_�G� �� 
$WARN�M"`#!�!�p�@LI��f�NST� CO�R-�RFLTR^`�TRAT;PTb�>� $ACC�Q���N ��r$ORIأo"�RTlP_S�FgB�HGz0I���bT�1�I�ʐT���K|�� x i#�
Qnr�HDR�2J(; �3I�2D�3D� �F�5D�6D�7D�8�D�9�" ��CO�D <F ����8�#�܀O_M��� t 	PE�q0�1NG�1iBA � Q���q��!�Qp �0=q�0I�P�PJ�Y��G�S��p@m �RC �����"J��S_R��gC��J��L��ļJVep�%C�`X���p0�T�A�zOF� 0  @�F RO��&9�6�IyT3c9�NOM_y<V�lS 0$��D �0��A�B�'&�EX��B0��Px���
$TF�lE0��D3N�TO�Sr3U8P+� -0�P_H�j 1�E{� %�Y#&�d%(���1�$�DBGDmE}!_p$���PU��1a2)��I"��AX�Ae$]ewTAI�SBUFiv�XY�/ � �k�f�PI�$*��P��M��M��^�z��F��SIMQ� ��$KEE:�PAT0�����N#��Y"�4$�L64FIXb/��⥟TC_��b� ���c��CI�Ύ�PCHOP��ADD��������I"m0p�3�_��!f�� �n!
��a��W���d"m#�MC�� �0yJBE�ͤz��l��+�i�  �N���� ��pCH� EMP�$G�����p�_�lS��1_FPpm��@��SPE���lPn�������� V`�q<r�A��JR�~<rSEGFRA���3 �R�0T_LI9N{sMPVFs!��'�_�"�#m�"� �R�B�y0z� D )���`�����2 �f�)P���Ţq�f�SIZc���T���3�RSINF��G�R �@e3 e��> L�8з�CRC(�AcCCn��3 ���*���1Ma����D��D&�e#
)C+e`TAM ^�&��T(EVT&i�Fj!_
F��N�&�@f�`��((������'���j1���A! 1�>p��-�RGB��"��FB ׂ��De�RN��LEWر�Q����/�. x�|�Xs"� ���Ư�5b�#�R� HwANC�$LG~���!�QU�y�gp��6�A:`� a�c�R?2 �3`p0��3\��8RAnS��3AZ��7HP ��O��FCTC�Y07�F�)����R�ADI�KO�H@�@�o� �D~�.��6�S�p����qMPW*���M�4AES��l#��g����4#  z�I+$�CSX���H���$*�?p�s��T��B�C�0N�p�I�MG_HEIGH�mqrSWIDK��V�T��M��pF_Ap {��B`EXP�A�4��U�CU7�]�U�%�% $_�TIT&���r�s�p��LE:RZ_% {�&*��{� ��A~�NOwPAD	q?W�i?�,����D�DBPX�WO�&�'��$sSK���r  8�`�T�0TRL%�( �,�A!���@��r�DJ��LAY_C�AL�q	��`�@�gP�L	�G�SERVEADW�wb�w��'���	���9��0���Ȉ`AA%�)�b��PR~� 
��D"����%�* _����$�$"��eLoy+|"ф���&�,�"���PC�%�-�"Ѩ�PE3NE���!.�"��HOqRE}��r/�H�0C�� *$L2�+$os��+@�C�T ��O�0_D�A��RO�����䤍�|�RIGGE<�PAUS��V�ETURN���M[R_�TU>���a�EWMF��GNsAL����$LA-���n�,$P��g-$P\@!�.��b��C!�!��DO�` ��\�H��b�GO�_AWAY8�MO�D�0�B,�DC�SrpEVIm� �0 P $іR�B�
�PI���S{PO��I_BYT2�����TXw�L$�1� H� 7��Ф�TO3FB��FEl�������w�CU2�D1O����0MC��N����7�`����Hy@W����� �w�ELEGR3 T����cCGINKh�����U퐍L��HA��}y$��} <w�ܕ���4 ��`MD=L�� 23��(�!O��^����C�2����J]�}O�m�}�2�U�r�h�������	Ĕ����`W��45� $]��0�PcC��PZ��Pa5бw��ϲ��̵IDJ�˶�br˶W ���NTV��вVE��(РW�D�	2W��J�&���p�SAFE)���_S}V�BEXCLU�a:��>2ONL����Y6��3x@�Qw�I_�V�@�PPLY_`���� Ƕ��_M�"}��VRFY_�c��MS3�PO��x@!�"�@1~S4�^�O����8���@� 6��`�TA_ ���� �  |��SG�  �7 ��CUR�π�}S��tpUQO�R�EV�ٯҦ�jPUN��p��ԥ��Ё������0���ѧ@��� ���PаI�r8� @� F���T�OT�At<�At'qAt�^� `+�M��N}I�r9 L �`���Aʱ��DA=Y	�LOAD��6t4v�Bs5w�EF�P$�JX�:�' SO�����P��`_RTR]QX�; D�!O��RQ{�������:| C7 � �qA;`���< 0��Z��p�Z�>��6DU�5��bCA�� 3=9�[`NSk���ID� PW93U�����V��V_U��< �DIAGr��u>8 *$V��T%ep
Dp}R�r��{V2`7��SWB�� u���R ��;�� �3OH�r�PP2a}IR�Q}B���m�`����|	�BA�����D@������=���CY �RQDMW�MS� AZ`xw0{LIFE�`�/Hq��NB�K@��@��!����C�@+f�NЀY0�QgFLA�4��OV�@�W.`��SUPPIO�`�A���`_���z_X�C�a���Z�W��A��B���CT%U? `>��CACHE�'C"�ۣ�կ���� SUFFI�ϰ�`%a�6t��Bs6>q ���DMSW%U@ �8��KEYIMAG��TMF�C�!с޻&INPU}R ;��G�VIEL �1wA �BGL/�����?� 	
dnpfPcBMP�!g1CIN^�Tb��	UBv�JB���d��O#QT�3��S��Uu59d�;��OF��H���C �Va!gOTF���ץ1�D[�P_GAI�Q���@�@̒��NI_�0C���5��\�6�PTIC��O�P E���"��}1�A{�P�CF�@INy��P[EA�q�@!� ��A|$P�3D  P�*�6D�7I�8T�=ĹRv�=�AVE�FF�BP�c�C���3AW_�@<���E����;DO<4SLO���1TERCE/���D1L/`�J3UFU'RQ��E�e{0�P�E}1�D��B�FE��3N� �3qPQ;`�5�R�6�R^�5�G�FF� 8䠣�$2��G �1�0���1F ����0�3�0 ��AbyB��cCARRg#i0�9T$ <2%cyftqcRD_4�06FSN�p���T� �FSY��D�I"e�C��A�DĔ�dEG�R�F 	cu0��Hb�C9�0�ǰY���1�@3�GG  mq61��I�  { _��3]6�0�s�1�s<�1�r ��D Ц$�J�z�STp@!�r)��tk��tv��t<���pEMAI����/1��� �@AUL��K�")8}1COU�dP�!�pT!���L�,�@�M�SU��IATh�RZ�U'}�N��NF SUBRT��C�p�1�*rw�SAV~�@� ES��m�����r��P��M�ORDM��p_RPd���ډOTT���A�3P�60���s��AX��,��X8RP�R�YN_�>�!Mb��6�௕�G3���@IF� p����b=�N� ��05��r�C_RO�IK�"���Ҟ���@R�!���8��DSIP�&��PA��I(v����ß���U���D��M�pIP0Á���D  ڔTHRE�S�`˕��TZۓH�S�bۓR`�E[@��V�����@�㑤P��NV��G����]�ؖRP	FB��d���@(��!#SCbRu��M-P���FBCMP�À�EiT�a��O�"FU�cDU'��QPPEP����CDљ[���-3\��� NOAUTO��P�$z���z�V��PSy�CR���yC�BE Dv����QH��в�� r�г���@N����S ��k���v��������!*��7��8��9��BT���1�1�1*�U17�1D�1Q�1^ʕ1k�2y�2��2��2*�27�2D�2�Q�2^�2k�3y�3R�3��3*�37�U3D�3Q�3^�3k��4y� �v�OU�T� ��R � �"@	WvPRuPLCWCAR+v�`����R𾠳$FACm�S�E��$PARM1��2m�"k���x����pA�Ph�EXT���!S <�)9I��g�0Rv��枵�\�FDRdTT @ ����E�-�BE�11(OV�M�4T�A\�TRO�V\�DT��|�MX���vP&�{���IN	D��:
���`E�PG3���� b1�`�DRI�@c�G�EAR�1IOQ�K�L��N�@:EFF�\�k�� ��Z_M�CM1�E�F�U�R5�U ,��V�?g �0@?� �Ð0�Ei@� G|�p��2� V�R�TP�$VAR�I�5����UP?2_ W *�?�cTDI�iA>�TV���  D�BACG�X T�p@�U��=0)$PROG�C%?����B�ICFI�� wYPa���!��FMR2>�Y ,�k� �B-�Mp�1�8J\s�}0p�L�_���A�C@IT_[U�C_�LM��(DGC�LF����DYt(L�D���5����������uZ�)� T�FS؀�t[� P�P�":2�$GEX_�!�(�!1'��נ���!3;56�9G���\ ���2��4l�ON����1�TL�1Q�GR��U���BKU�O1�� ��PO��9�0�$�W5�0M6`LOO���1SMw`E�� �����`_E �] {�����,PM�5^�6  O�ORIp�1_
G�SM_M	�0�`�5�wH�TA�/Ia�5 �U�P:P b� 9-��b]$�5v@�^��G{J� ELT�O�CUS�@ONFIG��A� c1aC�rD_$U+aא�$}��A�@P� OT��G��TAk�-�3SN;STv`PAT`�f`�RPTHJ(�N�Ep� ��W��BARTE` �E�p���r�AR[pRY��SHFTR��AQ>CX_SHOR1�K�J.F 9@$HG�Pa>!�.�OVR����PI�tP;$U�� M�AYLO0�!A��`� ��pQ]���]�ERV� �Q���Z���Gv`QR��0t;e��tRC����ASYMt����AWJ�G����E�?QkibQ�U�d@A�CU�q�P�YUP��Pġ�VO5R@M��?0�1 �c�r�2�6P�@!����q�%d �t��xLTOC�A��1i$OP@o"����2��pH�YO��Z�REbpRأ���)�K�ReipR�U�u}x[QDe$P�WR$ IM�ubR9_Xs8TVIS/@�bsH,r�B e� �$HC!�AD+DR�H�1GR/�$���v�R3�����f H��S��N��� \���\��\�*Â�N��U�p�HS[�M�N�!g `uB�trq�[�OL1���h���^��0ACR�O�p�AhqND_C�1�|�a�tšROU)P��!r_ÐI1�Uq"q1��6�2��<��� <�Q�=��<�*�<�7�66�AC��IO���D7���G�X�� �gh $� Pp_D��x�0�⣂PRM_+�� 
`�HTT�P_|�H#�i (��OBJE���t[$�LES���ְjN0���AB%_��T�3P�S�����DBGLV1�$K�RL�yHITCOiU@�1Gf�LOC�=O�TEMPt���0��zpv{pSS���G�HWe��A#�kW�}�`INCPU���pIO�e���r������*�@�IBGN�$l���� 'WAI�s�aP�����R���FW$ ېLO�m��s|���y�AN�A$Bo�����p��������RTN/`��CUF_DATAp�㖠����_MG�2(/ F�>�S(SE��r�N�8REC���N�b�<2�h�I� �m @� N�_h�Y8�3t���EXEwɒ�.Ф _�Xu�0�}n�$SCH�`�QP�R��FLGBvQ ��3�	/�oo�0����v ��OPÒ�1~�TRA�B��CS�D��9�pxw $C�CTA�\�'�IGN�MoO҈0�M~�Tֈ���v���vN_PCSqO�QUp��ECFBa ��Q���u��Ғ�	\r���L�������@DFpRs������SPT �<$���SEQ_� Z3NS��H�*�ɀ��rC�q�@Xl�SL� }Pr�Q �-@o�bc���0�se:!��IO�LN4q 8��R��$SL�$�INPUT_�I$�p��P- �����SL���!rr��#��0��ݐF_AS:�"s:$LO$� O��Р�r+�����P�HYP���^� 	 �8�UOR��#t ` J��(�%�s�%�|����pP�s������|������ �UJR��u � N���UJOG�G$D=I,�$J7�d+J8O	760I�AX>j7_LABQHpxZ �NAPHI� �QY�D� J7�J8�0_KEY�� �K)�L&�%v � �AVއP��CTReS�FL�AG:2��LG�$w �����Y3?LG_SIZJ��0`>� =A�=FDHI<S�1J;@= :tsC�� �A�pj�@�X_R��x�����5D�LNC
H2x����U01#��!BpU�)!(�L�2#("DAUN%EA`�)�Dtd"Z GHEr� ��M�BOO>Q�yt Bd��pIT�Ø${�e�#ү('SCR��`�D��[2�$�MARGI�D��,�X�ct2��M�S�0�L�W�$M�=$X�J{GMC7MNCH�&M�FN�F6Kl7q�j9UFx8�Px8n�x8�HL�9STPx:V`x8àx8� x8RS�9H�`�;U�C�T�3�bX�p7CIU䑌47 �R,6� +�2G\9lPPO�G�:�%�3�d2�OCG�{8���GUIj5I�3�B(3S 43Sh0l1�P�rC9���&�P�!N݁-�ANqAM�Qq�QVAI� ��CLEARfD�n�HId�~Sr�~RO��XO�WSI�W�XS��X8lҸ�i�i1��T�քn�DEV��	���!_BUFFqzj� �pT0R$I�EM����' 0(
bjqq{� �p���ˁIpOS1je2:je3ja �
b~Q	p| �! ߈�aZSq��{���IDXtAP�ƞ@z�jK�T���Re Y���a {$EvC{T�㐜v)v ��ch�} L�s������`�����w3��u�Kc~�#_ ~ �� +�#��!�sx�M�C" �! C�LDP��vUTRQLI� wT2 �y�t�� ���p͑�nQD���ڠL���t�ORG2 B!�'���������!���s͔� �����tE�t�SV�_PT�p��R�Ǆ>φRCLMC݄m����MISC�� d%!�aRQz����DSTB���` K��!X�AX�vR� [�t�EXCE�Sm �-�M���⡂��?�vT � �p/��㠃�M�_�I�����r����P�MK�� \��P�MBۢLI�CL�B� QUIR�E,CMO>�ON�D�EBU����ML���Ш��e�8H�Pށ���2�5Di $D�$xU�PyACKED�����DPxv��IN�b$q�_Q �pI�U�� �����/�	�=�U��4�T�I��MND:!SSb�#""$f��DC�6$IN]ю3'RSMD ���PN�r�BC���y�P{ST��� 4q�;��fRIl �e�e�ANG�bI�����AQ���;�$3ON,"�MFq T��i��00�uz� 3��SUP�� L��FX&�IGG�! � �ဃs��#�s6F�tR{�v��b������ȵ�����+�DAsTA���ETI8 �,�Bp�MH�b� �t?�MD?�In!) M���YӇ�U�H#�S�X�DIA�Y�AN�SWe�Y�Pa�AX�Dl#)H1�ŀ���� ��CUSVؖ��+�����LO�f �������G�����5����� � �t�MRR22��O� ��J!Á� d$CALI�Q��GrQD�2f`RsIN�0G�<$RR��SW0�����AB�CS�D_J2SE�e�I�L�_J3��
���1SPm I�P�����3���ѓ�I�B��J����āOa�IM��CSKP �z<�- kS<�Jm!��Q<�m�S�m�c��_cAZ˂	��ELa<���OCMP&�����1�� ���`1����� ��Z����OINTEVpSb����2I��Vp_NB���7�a'��3̒�A	DI����`�DH��6 ���Y`c$VQ঳�a$l1$ �!`��Q��-�2��H ��$BE���	�qA/CCEL����>� IRC_R-���ONT�a�c$P9S���rL  �!��s -!sPPACTH�	Z�Z3)����_ga���ʂr�C��� _MG�Q�$DD��"$FW5�1�������DE�PPA�BN1ROTSPEE�ka/�pc�ka�DEFۑ�)$OUSE_P�>SPC�@>SY
 � ʁ �aYN1�Ac�x&,��o�x!MOU�NG�tB�OLJ�$INC�� ���X��'3�Y�ENCSP��I��!�V�IN�bI`)52��c�VE� <H�*223_U>��^<3LOWL�Qz@���p�%\6D]@I�3�� �p�%�C' #6M3OS�P�MO���`�ʇPERCH  y3OVp t"�7�a�3 ��_2�������b%�$�P*�A)EL=T*��)�$5��_:ZFu6T3RK�4�bAY��C ܑ�A)�E�C!��`��RTI���"�`MOM�BX�ܒc���G���D��C\jb� DU�2��S_BCKLSH_C)U� �6 �0�#��:T�"EZ�!e�CLAL2`"2���@��`wUCHK�p�eSN� RTY���5�$�U�0�_�c�4_U�M���YC�S�SC�L�T# LMT��_ALg����T�gE m !`k�Pe��0Q0�!&@bd�8PC�1�8!H�pl���UC뀎rsXT� �CN__�1N���f�SF��9Vb""�7��a)un�hCAT�^SHo� _���&U�Q6��*�����PA�T�"_	P�U�C_�p�P�F�00�q�C�t�UJG����̧sJ0OG�g�BTORQUT ��3�I�`/��2�A��_W�E �D��7��6��6�UI>�IL�I�F9�`)��#�VC� 0R�䒬�1����Əc���JRK�����~��DBL_SM�!:5BM��_DL�5BGRV=�6��6����H_���]d�CcOSq��@q�LN�� ������� �� ��h�Қ�����Z���6�cMY���}�TH���1�THET0e5N�K23�[����C�B`�CB�CT�ASƱ��h������`��SB���k�GTSE�#!C�� ���|s��<�ϓ$DU�P>G��D��!���3��AQ���&�$NEB��I���#���L$~ O�A�S�|���c�n�n�LP!Hq�Z�45Z�S��ͳ ��ͳϕZ�ޖ������~ V��V��� ��V�źVһV�V�V*��V
�V�H������µ�:q��һH�H��H��H
�H�OJ��O��OIٴ�OźUOһO�O�O��O
�O��FZ���������ԑ�SPBAL�ANCE�~aLE6ȠH_S�SP���4���4�ϖPFUL�C8�_�G�_�ϕ!
1=���UTO_�P�u�T1T2���2N �Quc���O�Aa�?�(0��ATK@O���>'�INSEGu~1�REVB�~01DI�FtEF	1�+�r1�g@OB!�gQ@��G�2����Q�LCHgWAR
"g"AB�q~�E$MECH��� ��!��VAX�AP�Ed��u�� � 
p����5ROB�0�CR)���b d��MSK_���� P ��_R R ���+:!vD1r/0�-"+ ,3ET+ �IN���MTCOM�_C��� �  ��3� !$NO�RE3��OPW�O��� �, �k SBU��QOQP� �T�
U��=PRUNq�P�AR D�����0_�OU�!�S�AB��"$ IMAG�VQ( B�P�IM�� BIN'�BRGOVRD<��	@BP!Ap!_��0q��R�`RB�`���[aMC_EDTU_� K`Nl�M��JaPMY19Ia�|�nSL6�" �� x $OVS�L��SDI0DEAX�c&�cKA "V�!$N'!�5 %#:'�5(��Q ��_8� �" � @�pl"P���2� �2
&_��x�'�!�! !��0��ECT�  � �H(��PATUS�P{@CD�ZDXN�&BTM�'�!I	��4Ia�#�" � �D( E"�"Z�E<4��!FILEJ@gP�!EXE� �Q�72�K24t#�{ ) � UoPDATZ1$T�HXNDP�������9��PG��UB�!���!�!~�#JMPWAI'p�P*#�5LO`�F��p�!�RCVFAIL_C�A��1R�@� �V�a�d��<E��R_PL�#DBsTB�q�UBWD.F2� U�P/EIGI��TNL#p0D�B�RT�� ERVE��c�D�bd�1DE�FSP�P � L( ���@``�qp�C�UNI"7�@�1RXR0!�.�_L�P�!? ��Pr !�� 0�q�!] A�TA$�uNP�KE�T$R#�BUtPI�PB!� h�ARSIZEp@E0�GQ�RS� OR�#F�ORMAT��uDC�O�Q�EM��̟TSUX� :" �,�PLIpB!��  $| P_�SWIp�d"h����U@p@AL_ W� $�AAVB�ꅠCVD	$E6Z1�`C_zA� � � Q��VaJ3��V80R�TIA4hi5hi6~VMOMENTtc��c�c�c�c| B @A�Dtc�f�c�f�cPU��NR�d�e�c�e�b� ��S�P H$PIQ��6� H�Z�l�~���!ڦ������� ��GQ�&SPEED�G�R�tE �D�v�DE�,@�v���x��y�ESAM�#��F��wL�EMOV_AXI�!�z�@�%���7�z��@1d
��2dR	 md��	`a Б�INڌ	`/� ���؄B�#���#�C�GAMM��A��Rn��GET�rFIMS��PDcd
��LIB�R�1�BI�@bS$HI�0_^� f���E`ŘA���ӖLW�� ����$�Ӗ?b���@aCfEq�|� � $PDCK����_.��PdւSiaɅ���c����f��c �$I� R��DW��1"D��LEa�q�!��?hᠣVpMSWFuL1DM`SCR�8�6�37+�U��q� ��S]�p��P��URB���GR���S_SAVEc_D����3NOC`C�!�2Dd����Sj<v 幾Uy�mp����p�W�v<Ƚ�.aO�AA ��񊅰���e�x� �vv��ǜ�ZÌ��1� D�QMu� 7� ��YL5s~� ɇ��~�����NB�KA	���WѰ�(��A4��`�����M��FL�CLK�aD�Z^�1j�X�PM��~ � � $��ή$W�Є�NG 1]a��d��#d��*d ��1dV@��s���S��J	`XPO+caZ&�8�P@t� p�| ��Uv�����,�t;�Ca_�� |� Si���i��c��c��mj	���jE@��f S���y��f ^`���P�Q�PM4 Q}UP� � 88PqQ�𽡤QTH� sHO��HYS�P3ES����UEr��hP��� � @6B;Q#��#��_� 0'Ѵt���EN/	PBG_@B�[mB?�H#*#Jہ��I��pEW �vGTF�-b"�PO�4��   �𮗫"UyN� N� p{ �rp� PD�E���-3�BROGRA��!�264M ��I�Th@�{ INFO�� � ����	�� (àSLEQ�v6�u$6�{ �D�0p������Ov����#���E��NU��A�UT���COPY����0��qʰM��N8��^�PRU����} gQRGADJv!e�wRX'��B$P(&3�&W(P(��$�s	 �3EXF@Y�C��	 !NS��T� �4ALG�Ok�.`NYQ_FREQ��U �w�!�T�LAhC�!��b.���5CRE�0��l�I�FQq�NAT�%��$_GhCSTAT�@4��M@R���31�	���Q31��|$ELE�0 �Nb�SEASIr1���"� a2�1���6BƀIa��"�q��M���2AB$�Q/`E� �pVU1�6�BAS9b�5����U8�@� ��$�1F��|$��� X ��2 2�  	����QFBPGQ|�r��eE|F �|$�PFe1�=GRI�D��SB|P�wTY�s3��ŀO �1Q�m�� _4!E �BwsRO$��$� ���;LI:�PORAS�C\'v�BSRV0)T6VDI�PT_�p6P�HT��RW�pRW4PY5�PY6PY7PY84QO��PFs�e1�� ?$VALU�3��̅4��	��Q�$��| n5	��C
1���0AN���R1�Rp�!��TOTA�LQ���7cPW�#I|�AMdREGENKj`b4�X!G�s�&��f�m�TRC�rKa_S���g``�3V'����c>�1E:3�@��ܚcV_H�@DA8}��`pS_YƱ�ڻ&Se�AR}�2��>@CONFIG_CSE��`RJ5_� ���Q�E� 4�{�O�v�k�F�PSܢ�F�f�C_YF��m���L�����(cMϰ���q�rd^⃁z��DEհ�2�KEEP_HNADD�q!��0�	CO�0+��A�r%�,�Of�
���q�,��1��,�REMC�@+����Bh����U4�e+�HPWD  �q��SBM!�0�uB� ,?F1L�з���YN�p�M:�C���pQ�Er�� �l0DB�M�TRI�DA,�Bx� 0�K�TCLA�����U AYNSP��֡SEAꠁ�GK_P�Tn���B���RGIn�QSOL!UK ��P��)a&�$SC`0D�#ے�ALI�r���S��B#U�A}��A����� ���w1�_8�P�H�TIC[��`�p[�REVI�o��OLP���p�F�K��_F�SSEG�Q���b� ��ITc3� �l0CP��{TU� MSEC��MN���̢������`�0�G����0O��1�$N�̡_�e�$�PA� j�P�vO�iP��MLr P�� .~� { S|е��e1��  $OW-����G����p@���Hp2C�ĹAü(�!ߤX�AX�Q��A7HI��6���ٔ�2��Ϛ���B�V�EP���P �`Q���H�ߢ�r��V�t��`a�B^"�$4:�Q������p�MĢ�y�O��l""�SM�H��<�M=�2�� �L`UP_�DLY��ÆDE#LAk�>a2Yߔ���  <�QSKI�'�� �P��OF��NT\P�B��P�� ���`
��P���a�� v��l���vP�ڃP��@�P�ڝP�ڪP��9���J2#����yrEX@T�#z����z��.@�z������RDCa�� �s ��0TORq���	��!�����SD�RG��H��k���G�g��eER�qUBS�PC�G�z�?2T�H2N�!D�#�1�� ���@��11�� l�p2�F1�7��Ta��� O ѯ%��� �����SDx��VAHOME��g0]�2e��k�}���������� �]�3e������0B.�]�4e��ew����� �]�5e����*<P]�6e��_q����� �]�7e���� //$/6/W `]�8e��Y/�k/}/�/�/�/ X�]�Sπf��  ��AX^�u`� i]�ET�ypa��m2.fk3IO�pr�:I0�� �]��POW�� � qU0K��� �]��(d ���2$D}SаIGNAL#g�f�CJ�1 ��R�S232q5� ����%8��ICE`t����³��ITq�&aOPBIT"cF7LOWCpTR003bZ��UXsCU+�M�S�UXTđ��I��FcAC1Dų%@ A;CHQ� @{p�p���C�$�`�`O1M,p_���ETޠ�s�UPD�pA3�  ��	@P�@�Q��+ !�(s�A����x�)��.�ERIOc�E�PT:p3T�2_��0�Q/PDAMVWR���/�9D��qV��6FR�IEND(�@�UF�i��t�P���UMYH��p@���GTH_VTE�TIR���R��P�XUFINV�_��ѥ�WAITI���WX���Y7fG27WG1��@1S�Qbbgpp_�RE�O_@t��s�Q�`��[PC�C�u��_TC3��Ķp��eX�GˀŲtq��@&Q/A�r�jQX�E8V��Ea��������D�X s�ML����`��SX��]E�#T�CG3�WCPgw�s�|tD�LOCK�kuvӮ�V��q�ta�	$�f[���pkQe�qY�1}XlP2o[2�{3o[3}Z�y'�~Y�yC�`6.�s.�r$VV�J�V8eVl�� �a�b!�غ��F�sρ ��fqB���`�R�ɠ��E�$߂�S�@0a�Tu���PR����uj�Sl�G��f3�B��� ����%s[��w���[���p�@|`�@Ҳ�
\��BS�1� ؚ�R_6�oQ����`RUN��AXSA�`A�PL�QV⮒THb�J���6�aq�TF"�NT���IF_CHeS��~�qU��6��G1��0�t��� 6�_JF?�sPR�`���RTC�� ���GROLf�A�MBVq̐Cr�̃��`UI#���BU)cRSM}��a`r��_W�P�TBC_-P�PCM��D��ЖLDR��ރ�A��@���c�IT�" �4���TA���# s���|� �ҙ���� ���� ���2�  2� ��S��g��	| �Vд�}�I�t�ˀN~�TOT��~�D�>��JOGLIzC
`'E_P��qBO��}�����`�FK��_MI�R��Ѵ{`M>r�A	P]q��E)P�ҔJ��SYS�˂J�PG'�BRK�bѕߐ��I"1  N�pSY�Ā�x�D�A~��BS�O�}��0N��DU�MMY15U�$�SVVpDE_OP�oCSFSPD_O�VRU��� LDL��óOR��� NPb��Fߑ�Ʈ�OV��CSFڟ��.�F ��́ճc8ؿQ˂LC�HDLz�RECOQV��[P��W�PM���vձ�ROoC����_� ��� @�&`V�ER��$OFS2&`C;��SWD��r�`����Rū�TR�1�W1FpE_FDO�ƃ�Ӡ��B��BL �����1K0%�V�A�B��@��b� �G�,�A�M*Ã�D�Z��t�_�M0�|B��3��T$SCA���DU����HBK�AЖ��IO�oU��1qPPA �����������2��?DVC_DB)c0�@ё�21���́H�1P���H�3P���ATIEOˀ�A{���UtS젆6CAB��nR�c@7p���`S��A��_�@~ЖSUBCPU�2��Scp�0�B��@s�j�B��2��$HW_C_ dЧs5�s�Ata���$UNI�Tb�\ U ATT�RI�i��CYC=LϳNECA�����FLTR_2_FAI��8���6��Pǻ���_SCT�cF�_UF__�q
FqS�1:�ZCHA�Q��)9�qB(RSD����2x�ޣ�1�0_T�W�PRO����g@E%M*0_��V�Tq�� z��DI�PҔRAILAC4>��bMg�LOu��S��9�R܀��䁟���+PR2�S�a�p!�C$�$@	��FUN9C���RIN�`Ԥ��'$fARA8 �b ���P#X0��P#WAR/���BL�af'�$aAz+v}(v(DA`�0Q!�(�#z%LD�@���q�#��Z!ہ�#TaI�5y���$�@gRIA�A�2AF��P;A.3��45�p�r�@�MOI` ��D�F_�P7��Ac�LM���FA�PHRDYJTORG͢��fS� >�5MULSE�P�T���J��J�������FAN_AL�MLVV�AWRN	EHARDpP�E��Y"2$SHADOWl��/�?Bc�@w@du�:�_m�ЖAU�`��:�|@O_SBR &�E���JU &�/!�C_MPINF��k��D�!�CREGpU�8�л�i�� �`�Q�$;Q$Za�e�O�j��� ���EG�~���*QAR�����2�q7W� �,�AXE��ROB ��������R�_�]w�CSY_�dQU��VS�W�WRI�P=V5 ST�R����T���EWH8�FT�qkB�`B�P���V,�����OTOr�A8���ARY��`3b���B�ƱFI5�ܳ$��Kq1��Sa%]�_�S��EU3��zbXYZ'B�j5N�fOFF��RbzbJnh7`B��"�d0��V�  �cFI� �g�q��«�"��_J0��6���y�$a@d2k6��qTB)q�22arC� �DU��DV]7�TUR@X
3��uAa�BX�P��IwFLg�Tд�7P�p�e�Z��û� 1�8�K��MДDV����ORQy��V#�W3I��2�+�s0�h�tà�Tz�OVE����M� *��C��S�� 
R��6@��*A��W �� <�! �50�����݀ Q�*�������'�S'�L��ER��Z!	�!E�PD��e�A����eH%t?g�!���!AX��6��!Ua ���˙�1˙�`ʚ�` ʚZpʚ�pʚ��ʚ�ʚ1_�ʖ�0Ǚ�0י �0癮0���0��0� �0'��07��0G�d�X�oDEBU-$(!`4C����vbAB������~�V��, 
#�Y�?�K�OW�#a W��aW��aW�ZqW��q W���W��:4fp42��.�cLAB�bI�) �6�GRO� Ir-L��B_�L��T���`��@ �4�J�0�A<�AND���Z���e]�Ay� ���@~a�ȳ!��ȡ ~`NT@=!��SERVE��P�� $0 T Ae�!��PO��K@��-`���0��_MRAQ�/ d � T��e��ERRr2�00TY2�I��V�`��7�'TOQ����LhP���RJ� ���D@Q � p 4�����_V1f����Ԥ
��2��2���D@�pq�H����$W� ��� q�VQ��@�$���d0i�x��O�C�!P�  ��COUNT�Q ���SHELL_�CFGQ� }5!pB_BASVC7RSR�AB� E~SSW�!h�1��U%g�2��3��4��U5��6��7��8��[�ROO�0��Y`}`3NLQlsAB�úni�ACK4�IN�T� ���0a@�0��_PU�0@�OU�3Ps l��I�����TPFWD_KcAR<ї0�RE���0PO`�! QUE�r�t��� �r.@_AI @7�H�{`�D��EzbSEM?Ox0)66�TY*�SO��)�DI6�s ����b1�_TM��'NRQ�g{`E� (�$K�EYSWITCH����I��HEupB�EAT�qE:PLQE;��U��F�����SNDO_HOuM20O<#REFe��PR�a���Q�P7�C"� O�1�v�O �;r<K@0IOCMgt���a� \G�HK�Q� Dxat�RESUUB��M�"��w�wsFORCx�#\�|G�OM;P G� @�*3~@U�SEP9P1�$9P3�}4� ��S��HDDNP� ��BLOB  ��pPNPX_AS�P�� 0v�ADD|�GA$SIZVA�$VA:���0TKIP�'#�A�?� � $c�( H�`bRS��"QC7О�&FRIFHB�S����� NFjODBU�P���%�#�)>�� ��Si�P�� x��SIT�TqE�sX��sSGL#1	Tab�p&��<3íP�$0STMT�qU3P�&P�VBW��%4SH�OW]5�ASVDT�U�� ��A00~Ħ2��7��7P��7 �75�96�9U7�98�99�9A�9 \P�7��7ӱ�6�P�7��C�3W�pH�91�91��91�91�91�91�I1I1 I1-I1�:I1GI1TI1aI1
nI2�92�9`@X�9 �`@X�9Yp@XI�p@X� I2-I2:I2GI2
TI2aI2nI^�h�9U3�93�93�93�9U3�93I3I3 IU3-I3:I3GI3TIU3aI3nI4�94�9U4�94�94�94�9U4�94I4I4 IU4-I4:I4GI4TIU4aI4nI5�95�9U5�95�95�95�9U5�95I5I5 IU5-I5:I5GI5TIU5aI5nI6�y6�9U6�96�96�96�9U6�96I6I6 IU6-I6:I6GI6TIU6aI6nI7�y7�9U7�97�97�97�9U7�97I7I7 IU7-I7:I7'�7TIu7aI7nD d�0]P� UPD���"�+���
h�0GUN{_C��� `�ng�PUT'�IN\����<AX|�GO��U
GI��IO�_SCAw�0YS�LOP�� �  E%�"#��':'� d�� @ʤ	�P�� �R��=F��ID_Lj+��HI&�I���LE1_g�V���$	 v��SA��� h�~��E_BLCK�����M1��D_CPU���F ��: &�Y�k�4x���b�R ��g
PW"��� 	�LA�2S�����RJ�FLO5��5��đ 8�V��V����TBC#�C!��X -$}�LE�N��$}�D�RA4��d!$��W_��&�)1}�C�2��M�b�h��� 3�II� ]ю��TOR��}��Dx����� LACEG���}������ _MA�+ �J� �J�TCVQ�r� �TssڒՈ�@���� ���JF�&�$M�ԙ�J���0R��� ���2/ `~0���ӱ�JK(�CVK:�$B�3,�J0O�>�JJF�JJN�AAL>�t�F�t�n�4o�5��NA1�ܥ�d�N�y�L��n{� Xx�CF/!��T�v�M?1�"B>�NFLIC�# REQUIRE�EBUOy���$Tx�2�6�z� �x��. �3� \rA�PPR,�C��{�
���ENs�CLOS� ��S_M� $ ����
�$��A?  ������  �����%��������s�VM_WRK 2 ��� ?0  �5��B)L L	#�`������q���_��n�+5UXѠ;M _�������/B/T/7I�)$ORk}�5/�/ �?�/-?;?1/r?��?g/y/�9DYN_ �/�/�/e?O�/6O? O?]OkOa?�O�O�K���BSPOSU� 1���� <�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
���B~�N�gLMT�����C7  �1�IN:�L��0�PRE_EXEb]���l�.�AT}���J����LARMRECOV ���l��DLMDG � "�LM_�IF ��d �*�<�N�`�n����𣯵�ǯح, 
��O���FNGTOL�  �K�@A  1 4�F���PP���N ?�������Hand�lingTool� �� 
V8.?20P/A2E���x.p
881�50���80��3�348966��x?is
91����pra����rod?7DE3����pc 	F�.�014i�Y p�FRL�ld�32���V9�X��TIV}�l��J�i�UTO�� ��h�P_CHGAPON=���������L�1	� ���������I��Un� 1  \�
���>j��4�����VIQ�c߽߇���{�� �{�Ʋ�HG�����HTTHKY�ߚ߬� ����6�H�Z�l�~�� ����������� � 2�D�V�h�z������� 
������.@ Rdv���� ��*<N` r���/��� //&/8/J/\/n/�/ �/�/�/�/�/�/
?? "?4?F?X?j?|?�?�? �?�?�?�?OOO0O BOTOfOxO�O�O�O�O �O�O___,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o �$6HZlu*�T�O�uχ�DO_C�LEAN��(��sN/M  #��9��K�]�o����_DS�PDRYR�'�H	I���@(���� %�7�I�[�m������8��ǟ$�MAXZ��t�q�q���X�t����|��i�PLUGG����w�Å�PRC��B��ϋޏП?�OxD���(�SEGF��K�������'�����%�7�o���LAP ̏߮�Ӌ�������ӿ ���	��-�?�Q�c�>��TOTAL�0����USENU̠��� �x���r*�RG�_STRING �1��
��M��Se�
��_�ITEM1�  ne��0�B�T�f�x� �ߜ߮������������,�>�P�b�t��I/O SIGN�AL��Try�out Mode��Inp��Simulated��Out��O�VERRɀ = �100�In �cycl���P�rog Abor������Stat�us�	Hear�tbeat�M?H FaulD�M�AlerW���u��� ������������ �s���q� hz������ �
.@Rdvp���.WOR�� ���X�//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b>PO��8�0�q? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O��O�O�O_�2DEV �>,P�?_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�oPALTD�a� �o�o
.@Rd v����������*�<��oGRI ���t��oN������� ҏ�����,�>�P� b�t���������Ο��b���RD����@� R�d�v���������Я �����*�<�N�`�xr����PREG�n ��0��������,� >�P�b�tφϘϪϼπ��������(ߊ���$ARG_�D �?	���k���  w	$��	[��]�����^�SB�N_CONFIG� kۊ���C�II_SAVE � ������^�TC�ELLSETUP� j�%  OM�E_IO���%MOV_H!�4�:��REP���X�UT�OBACK�
���FRA:\Ϊ� �調'`r#������ ����x�15/�12/03 07�:34:46����ت�B�T���x��������������"�����Pbt�� �5���( :�^p���� C�� //$/6/H/�'��  ��_��_�\ATBCKCT�L.TMP DATE.D�l�/�/�/\�/��INI�`���֞�MESSAG����!��s�����1ODE_D&����-(1�O.P0> 4PAUS��1!�k� (�7�?I���I?2������n��g"6�+��)�sB��諾9����? I�?O  (On�(O:K$OZO�HO~OlO�O�Ic4m0TSK  s=�1�M>�/OUPDT'0�'sdP5XIS��?UNT 1k���� � 	�@�M�D8)� ����nKS���A�O�GQ��� -e� 0��M (~ �h ��b^�_�_�GQ�j��$��|7 �g8�ݢ 8OM �_�׭_�_oo=o(o Moso^o�o�o�o�o�o �o�o 9$]H �l������ �#��G�2�k�V�h������ŏ���T�)QM[ET�15]Pޏ 7�ڏ[�F��j����� ��ٟğ���!��E����SCRDCFG� 1k�u���X @� ����ȯگ�����"� ��E�W�i�{�����
� ÿ.������/�A�0SϾ�YԤ�GR.PPXQ?}�j NAN�j�s	��z�_ED� �1t�� 
 ��%-p EDT-�k�b���߻�� E@�-����/��ґ�?���.�ߗ�0023  �����2H� ���$߾  9۹�$�k�}��/���!3\��ߩ��?�;R<؀����7�I�~�1�x�4 (�F����d���Q��� ����9���5��d� A���������w��6�0T����T��C���7 ��� ��� /gy/���8X/��/����/�/3/E/�/�i/��9$?�/q?�/� ��M?�?�/?�?5?��CR���<ONO�O��O�?�?qO�?}���N�O_DEL�ϛ�GE_UNUSE�����LAL_OUT7 ��  gҜ��WD_ABORT�
_{�CPITR_R_TN  /����~CPNONSTO���nT ���$CE_OPTIOkX��ƣPRIA�_I	PnU�P���PFn�+[ڳ/���Q_PARAM�GP 1+[�^g�Qocouo4k�C�  �n��`���`��`��`Ș`Ҫ�`ܘ`�`�`��  D�`�`*�`�`�d�`�m��a	��bD"p/��`;pH�`Tpa��`mpz�`�@ {D�p�� D�`/�?��o>ogy���n|�`��`��`��� C��p��p���p��p��`��`���`��`Ř`ʼpЪ�pּpܼp�p��`�����|; Mv���������� 1��ŏ׏���I�[� m����������-�?� Q�����	��i��P�HE�@ONFIG�K_��G_PRI ;1+[ t�� د���� �2�D�V����KPAUSPO�S 1���S ,]E������ƿ��� Կ� �
�D�.�T�z�@dϞψϮ���j�O�Q��_��QO_M�ORGRP 2�l ���Bs7y=r�:� 	 :� R�@�v�dߚ߈�k��� ����������2��� h�V��z��:�L�� �����
�@�.��c"�!݋���?o�o�H�`��0K���1r� ���������������P�P��+U��` Ua�- ��k}��:
\��	�0P�N@f��5g�`�53DB���+YI�2)cpmidbg[�@�m:�  +�	��UApG�k�`���pI��E���`;�a���-/�����`_��g/v/A/+~���fe/�/����/?ud1:��/?�7"DEF ���7)�!c�!buf.txt�?e?4 _L64�FIX , ��?�\�?�?�? �?&OOJO\O;O�O�O qO�O�O�O�O�O�O"_X4_F_~?MC�,P  d�_�_�UfS�t]��T�Ub_A�l�CpBp�:�B��wB���@B��LB�b��B�*'C<h���
;�D�6D��lD�9fD��	�DF=�D����mF6��F�7�F��+�F�DF�~�'F�&i�2���]<��YF	¬T_��;�I3`%�o�oL���o�lo~o�Y �oQ<u`� ,�����;��t�6g� =<�	J��������eأ��ӣ�x����`C><����<�p�  D��n��D�π��fE�πȏ  Ems�aT D�z��C  F�E��fE��fL���  >�33 ';��s�n����@s�5�@33�3�.�� A�=L��<#�
�2����/����� ��0�Q���Q��E��� �� H���1�9�J;#�H�2��Z��J� 9�Q�e�w��������� џ���B��f�=��� a�s���������ͯ� ���'�t�s�]��� ���ϥ���ɿۿ���5�#�v�2RSMO?FST 6>����9T1�PDE !=�pG����;�3�U�O�>T�EST02��R�7"r��|�| C�4�Pʀ��� ��J!�C�B���b��c�C�@i�-J:d[�
-�I_1�#7��-�T_00PRO/G %r�%v?���*�T_INUSER  ��(�C���KEY_TBL � ��(���@0�	
��� !"#$�%&'()*+,�-./01234�56789:;<=>?@ABC00�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~�����������������������������������������������������������������������������������������������������������������������������������������t���L�CK�����ST�AT`+�_AUT�O_DO�%�INDT_ENB�� ��П�T2<�-�STOP��wSXCh� 2$B�� 
 8
SO�NY XC-56�L輸�  �@���ʹt( ���OHR50�K��o�7��A�ff���//  �>/P/+/t/�/a/�/ �/�/�/�/�/?(??�L?^?�TRL��L�ETE� �	T_POPU��-��T_QUICKM�EN�4SCRE��0B��kcsc�4��0�9��c_�4UM��0U 1��  <K��ofOK�EO �O�O/ÁO�O�O�DF<���_�O_P_�LS�tart SM �Comm %IBSCMANS[_�NEndxV�@�U��0�_�]User �Cancel�RU?CANCAC� o��L
�RReset>�BURES oo 3_E_�oYoko�o�o�o��o�o�@Zang=e�GZG_-A�_ �ocuL^�� �����)� ���_��ZVAG_KO�NFIG.�RVW�)��=�O�؏s�-D�ateieL�%DATEI�1��� ��E��.�@���d�v��ß������П"bMa�cro Step� tt�PMSK_�}<��LWait� Monitor~3ashtpes0b y�؟꟯�����������VCYCLE PsOW�PPWD�x���� DOW��%	#�_MAIN�:�a�%Cb�NUAL��?�ZCD��&H��C�[�	���������?|(��$D7BCO� RI�Ќ5�#DBLOVRD��%�NUMLIM���d���DB�PXWORK 1'���ϩϻ���|����DBTB_1' (7�P�Q����s�DB_AWA�Y��GCP r��=��3�_ALU��?3��Y�5��$�_DBG 1)��g ,I���d����I�Ѝ� �вޟ��r�M� IS� B�@��	�ONT�IM�7�����)��
)���MOT�NEND���RECORD 1/��� �����G�O��B1��U�4������EX�ECUTING

 ��	����)��P������U�������Q�����/��������A���U7����a����@Rd���s��F���bU�B�2���z/���6~��|U�Ճ��X/=�������7��YU�}�� w�>/�P/�t/_/��8��P?'p_P'q`Э"�/�/�/�/c/?? ��E?��B�g?y?�?�? ?�?0?�?T?���/)O ;O�?_OJO�?�OOO �O�OtO�O_�O7_�O �Om___,_�_$_�_H_������_o*o �_No9oGo�oc?�o�o��o;o��TOLER7ENC@�Bȉ�N��L���CSS_�DEVICE 10���üƹW i{����������sLS 11 ,}��E�W�i�{��������Ï�PARAM� 2����TuTu~tRBT 24,|�8��<I�� �C�vd �*�����&��`T�h˴��?�g۶�p���  �\  '�g@��˴��A���F���p R���Ɏ��?�B���Ʌ�zɇă@��\�7��1���q@���Ɇc��Ɇ���Z�l� ��������Ưد�7��� �m��C�y��D�C�9��Ѱ�A���A�ff�AI��A;33�Ad �Ɍ��B�`pѐ��U�̱C>���BffB�;�-��B*갉�ֿ��ҿ�� }<�� �b� K�@ S�D�ɍ)�K�]��� E�sυϗϩϻ���� ��>��'�9�K�]�o� �ߓߥ����������� �#�p�G�Y���3� ���������*��N� 9�r���_ύ������ ������8!3 �Wi����� ��4jAS �w���c�/� 0/B/-/f/Q/�/u/�/ ������/��/�/>? ?'?t?K?]?o?�?�? �?�?�?�?(O�?O#O 5OGOYO�O}O�O�O�O �O�O$_�/H_3_l_W_ �_�_�_�_�_�_�/�O _2o�Oo-o?oQoco �o�o�o�o�o�o�o�o d;M�q� �������N� `��_��o�����̏�� ����&�o/�A�n� E�W���{������ß ՟"����X�/�A�S� ��w���֯������ ���T�+�=������ �����Ͽ��,�� P�b�=�k�}��ρϓ� �Ϸ����������^� 5�Gߔ�k�}ߏߡ߳� �������H��1�C� U�g�y���A�������  ��D�/�h�S����� yϧ�������� R);M_q� ����� %7�[m��� �/}�&//J/5/G/��/k/�/�/�/��$�DCS_CFG �5����!���d�MC:\� L%0?4d.CSV�/��#=��A K3CH
S0z��/#>^?�?.�  ���2�1��?�7� �`i�MU���(RC_�OUT 6�%��!��/�!_F�SI ?I �9#8AOSO eO�O�O�O�O�O�O�O �O__+_=_f_a_s_ �_�_�_�_�_�_�_o o>o9oKo]o�o�o�o �o�o�o�o�o# 5^Yk}��� �����6�1�C� U�~�y�����Ə��ӏ ��	��-�V�Q�c� u������������ �.�)�;�M�v�q��� ������˯ݯ��� %�N�I�[�m������� ��޿ٿ���&�!�3� E�n�i�{ύ϶ϱ��� ��������F�A�S� eߎ߉ߛ߭������� ����+�=�f�a�s� ������������ �>�9�K�]������� ����������# 5^Yk}��� ����61C U~y����� �/	//-/V/Q/c/ u/�/�/�/�/�/�/�/ ?.?)?;?M?v?q?�? �?�?�?�?�?OOO %ONOIO[OmO�O�O�O �O�O�O�O�O&_!_3_ E_n_i_{_�_�_�_�_ �_�_�_ooFoAoSo eo�o�o�o�o�o�o�o �o+=fas �������� �>�9�K�]������� ��Ώɏۏ���#� 5�^�Y�k�}������� ş�����6�1�C� U�~�y�����Ư��ӯ ��	��-�V�Q�c� u������������ �.�)�;�M�v�qσ� �ϾϹ�������� %�N�I�[�mߖߑߣ���$DCS_C_�FSO ?������ P �ߣ���� �"�4�]�X�j�|�� ������������5� 0�B�T�}�x������� ������,U Pbt����� ��-(:Lu p������/  //$/M/H/Z/l/�/ �/�/�/�/�/�/�/%?  ?2?D?m?h?z?�?�? �?�?�?�?�?
OOEO @OROdO�O�O�O�O�O��O�O�O__*_��C/_RPI����@_ �_�_�_X_��|_�_o�0o+o��SGN �7��r`�$���12-JU�N-24 17:�05   ���03-DEZ-1?5 07:3�aC`�Ab IY1=R�aH�ܻa�a�5n�`wasM� ��i�ZX�_�o���VERSION� jjV3�.3.2�lEFLOGIC 18�ٿ�  	Gh���Ny��]~0rPRO�G_ENB  �5dEs�`~sULSOE  cu�u0r_ACCLIM�v���s��sW?RSTJNT�wra3���0qMO�|�a��q/r�INIT c9=z���� �v�OPT_SL ?�	;��
 	�R575@ch�74jm�6n�7n�50���1��#tNy��*wK�TO  W��o�+v]V"�DEX�wdrb�C`)�PATH �AjjA\KJ�LTVL2113�50R01\ VL\ARG2\k��LY\���HCP�_CLNTID y?vEs Go� ǟ��IAG_G�RP 2>����R�ؑ 	 E�  F,D�E(p �D�5j��B�  =�+�B��C�f�T�CeEC��  C��C�G�SCEZXB��Gm:jf36�2 678901�2345��� � �  A����A�=qA��A�33A��z�A��A���RA���A��ߠ���5j֠Ba@o�  A�`Ap�,�B�A�C�C��`;B45l 5eW��Ba
բ���{�A�ߠ�ߠ�k�����G�Aď\�A��A�Q� 7�� �2�7�F�7�U�U�ߠχ��۠����������A�ffA�۠򠍿�����ÿտ[�_��Z��U�O�
AJ�ߠD۠>�8۠2�,O�&�8�J�\�V�_`��A[��Vk��P۠K
=AE��A?�8��A2��+�
�Ϸ��Ϩ����[��������x�q�j�c��\Q�AT۠L��1�C�U�g�y�[� ��v����Ѧ�-��=�G�I�>8Qy�U�-�8��bq��7�Ŭ}�-�@�;�\���p����m�@*�Ah�а��<��C�<�t�=��P=�hs=��ᗍP-�;��M
��<#�5lÐ��?+ƨC� � <(�U�b �4����A���Y�M�5iA@Ab?5� ���r������:� ������5YkM	?Tz�
�2-��J�G�-�2��C`�-�xC����}�
��/G�{CEY����ɦ4ZH������/��Ҧ�ED � E���D�����m�/  8����	����?R�?�Q��M@���$�?�$?�&L�?�C��*Du�Dd��p ���`�o/���/J�/�"5i�E)��>��\�O���d�/?}/�&??J?5?G?�?D` ����ϧ�?�?�>�?O OD�V��uWO�FO �O�O �rO�O�O�O�O _�O�O_d_v_T_�_ �_6_�_�_�_o�_*o <o�_Ho"o�o�oto�o �oVoHO:% ^I���i����J��>:��6�-� �og�Iw��������� ��	����?�Q��o x��������ҟ���� ���>�)�b�M�_� ���������/�� (�ϯL�7�p�[����� ����ȿ�ٿ���6� !�Zω?�?�?�ϴ��? �����+O=O/�Aߣo e�w��o��]߿��߯� ����+���O�a�?� ���!�k������� �'�����]�o�M�� ��/���g���G��� $J5n�W�� ��	��"Q�C U7�y���Ϗ�� ����-//(f/ Q/�/u/�/�/�/�/�/ �/�/,??P?;?t?_? �?�?�?�?���?O�? O:O%O^OIO�O�O�O qO�O�O�O�O_�O_ H_wωϛϐ_�_���_ �_��/o/ooSo eo��9o�o�o�o�o�o moo�o+=as �o�Y����� �'��K�]�;����� �C/�_ޏɏ��&� �J�y3�X���}��� ������-��1�/ U�g�y������I�ӯ �ǯ	��ŏB���f� Q���u��������Ͽ ��,��<�b�Mφ� qϪ��?�����ϙ�߀�:�%�^�p߂�LU��$DICT_CONFIG ?m���sVzP�egWS����S�TBF_TTS { LT
����VER��xQ�����MAURST�  LT�՜�M_SW_CF��@���ZP��OCoVIEW��A<�����ώ����� ����XR|��#�5�G� Y�k������������ ��x�1CUg y������ �-?Qcu ������/� )/;/M/_/q/�//�/��/�/�/�/?��PM�5�B<�xS��  ����;SCH �2H<�
�yQ�Schedul�e 1 LW ���R䑏9ZP?�?M�HA8�1�?L[=A�4>L�Ͳ2D �?�?�?O"O@OFOXO jO�O�O�O�O�O�O�O �O__0_B_`_f_x_ �_�_�_�_�_�_�_o�TJafeU4ueD5�9m*o �9Dzhg no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x�����@����ҏ�����5=`6�Jeb�t����� ����Ο���	H�V� �)�;�M��?�?���? u�;oMoo����ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ���_o�B�5�G� �7�I�[�m�ߑߣ� ������>����!�3� E�W�i�{������ ��:�����/�A�S� e�w�������S��# 5GYk}��� I����92�?`� r�c��T����ψ ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?��� �?����O(O:OLO ^OpO�O�O�O�O�O�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �&8J\ n�����@ R#�v��?�?�?H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d��?�o ���o�o�o֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tχϘϪϼ� ��������(�:�L� �o���������
�� .�@������ 3. ���6�� ��v�(�:�L�^�p��� ������������  $6HZl~�� ����� 2 D��p�x�ߦ�d߶ ����/"/4/F/ X/k/|/�/�/�/�/�/ �/�/??0?B?T?g? x?�?�?�?�?�?�?�? OO,O��P�O�O�O �O�O�O_ _f��b_ t_�_�����_��_z �V�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��PO8�tO�ODOv� ��������Џ��� �+�<�N�`�r����� ����̟ޟ���'� 8�J�\�n��������� ȯگ쯒O0_b�t��� ������ο�F_�_"�4�F���4��_�_�� �_��:�L�������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ��������^���4� F��V�h�z������� ��������.@ Rdv����� ��*<N` r�����R�� B/T/f/x/�/�/�/�/ �H�??&?�ϒ�c? ��T?�,���?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_>���_/ &/�o(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z���2/�/ ��&�8�J�\�n���@�/(?ԟ�`�5n� @?R?C�v?4��_�_�_ h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτ��_ ����ԏ揤����� ,�>�P�b�t߆ߘ߫� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�򏐟����* <N`��蟢��  �2�V�����ϖ� (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?�� ��x?�������?�?�? �?�?O"O4OFOXOkO |O�O�O�O�O�O�O�O __0_B_T_g_x_�_ �_�_�_�_�_�_oo ,o��p�o�o�o�o�o �o ��bt� �6����� z?�?V?��,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$��?PoX�to�oDo ������̯ޯ��� &�8�K�\�n������� ��ȿڿ����"�4� G�X�j�|ώϠϲ��� ������ߒo0�ߔ� �߸������� �F� B�T�f�������� Z�l�6���������� "�4�F�X�j�|����� ����������0 BTfx���� ��~�0�T�f�$� Vhz����� ��//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?r��BOTO fOxO�O�O�O�O&�h�__&_�z7���� �_��t_,��_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |����>�?� O&O�?6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v�������2O �O"�4�F�X�j�|��� ���O(_����`_r_ Cϖ_4����h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r���Я�� ���į����,�>� P�b�t����������� ����(:L^ p�������  $6HZl� ����//*/</N/�`/ƿϢ/�/�/@Z8 N_ �2�#?V�?���� ��H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ ���_����_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L��p/ԏ��� 
��.�@��/�/���� �� ??�6?ԟ�_�_ v_��,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� �_p�Xϔ���d��Ϩ� ����������&�8� K�\�n߀ߒߤ߶��� �������"�4�G�X� j�|���������� �����P��������� ������ f���BTf�*9�/��ҟ��� �Z�l�6��� 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/?~�0�8?T�f� $�v?�?�?�?�?�?�? �?OO+O<ONO`OrO �O�O�O�O�O�O�O_ _'_8_J_\_n_�_�_ �_�_�_�_�_r�bo to�o�o�o�o�o�o& h"4F���� t:?L??���� ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ^?o��4oFo o6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬ�Ro�o"� 4�F�X�j�|ߎߠ��H����� �10��k\�្� �ϟ��������"� �����j�5�G�Y��� }�������������B 1�Ugy� ���������Ͻ� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�߻�OO 1OCOUOgOyO�O�߻O �O�OYK�_o��R_ ��A_�_e_w_�_�_ �_�_�_*o�_ooro =oOoao�o�o�o�o �o�o�oJ'9� ]��?�?�?�?�?� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E��?�?�Oͯ߯ ���'�9�K��O{������a��$DPM�_SIM 2I����ʱt������C&]Y&Um� � 0�� DϨ�q���RC_CFG Jʵ�!�X� &]���ϸ������ ��5�6ᾰSBL_FAULT K���s�O�GPMSK � &Tb׾�TDI_AG Lʷհ�SQ��UD1�: 678901�2345��xz޻P �����1�C�U�g� y������������X	��Y�۽@��ORECP�ߪ�
�� ~�ܿ�ߴ���������  2DVhz��������9�K�U�MP_OPTIO1N|�[�TR��}�z_�1PMES;�J�UTY_TEM�P  È�33BȱЅ�A�o�UNIT|ׅ��Y�N_BRK Mlʹg�EDðZE|��'t�c�x�TA�T��EMGDI��[��NC#1Nʻ ��X/K/&^u�&[d���/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>COUOgOyO �I�!�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo �J<OFoXojo|o�O�o �o�o�o�o�o0 BTfx���� �����4o>�P� b�t��o������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �,��H�Z�l���|� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
�$�6�@� R�d�ϐ��ϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��.�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������&�0 BTf����� ���,>P bt������ �/(/:/L/^/x j/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?/O 2ODOVOp/�/�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_O O*o<oNo`o zO�o�o�o�o�o�o�o &8J\n� ������foo "�4�F�X�ro|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� j�t���������ί� ���(�:�L�^�p� ��������ʿܿ�� ��$�6�H�b�X�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ������ ���.�@� ��l�v������� ������*�<�N�`� r��������������� 
�&8Jd�n� ������� "4FXj|�� ����//0/ B/\f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �OO(O:OT/FOpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�?�_o o 2oLO^Ohozo�o�o�o �o�o�o�o
.@ Rdv����� �_�_��*�<�Vo`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟB����� "�4�N�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�F�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������ � �$�>�4�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
��H� Rdv����� ��*<N` r��������� //&/@J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?��?�?OO8/ BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�?�_ �_oo0O"oLo^opo �o�o�o�o�o�o�o  $6HZl~� ���_����(o :oD�V�h�z������� ԏ���
��.�@� R�d�v��������� �����2�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� �����Пڿ���� *�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮�ȿ �������"�,�>�P� b�t��������� ����(�:�L�^�p� �������߮�����  �6HZl~� ������  2DVhz����� �$ENETM�ODE 1O��  
����������RROR_PRO/G %�%��:/�G)%TABLE  �%�/�/�/��'"SEV_NU�M �  ���� !_AU�TO_ENB  q%�$_NO�!� P���"�  *�20�20�20�20� +10K?]?o?4HIS�#����;_ALM 1Q.� ���2<��+p?�?�?O"O4O�FOt?_OUT_P�UT 2R�= G @ٌ7���$_�".0  �01���J�TCP_VE/R !�!2/VO�$EXTLOG_7REQ�6�9S�SIZ_TSTK�;Y 5�RTOoL  ��Dz�2��A T_BW�D�@xP�&�Q-W_D�I�Q S�4�����VSTE�P�_�_��POP_�DO]_�FACTORY_TUN�7�d%iDR_GRP� 1T�  �d 	�O|o�m`��[���N�8�T&�hB�( ����fmc�o�m�d�A��?A� AM�ArxP��o�b��A���<A��@��R�o�oG2k�gA� ��AlA��N<@��>,@���P}��'��)l������������ӿ��|~P  <`�>�r���s=(��sz
? H C?q�u�Au${s�2_q�t E�  F�,DG�E(pO�D�E�4�D  E�Ўo�D��w�m��}C���N��B�ƈ����}@UUU��U�U��0�B��� �E�@���ԍOHcGP8��L�uS@�K�y�
ԍ?"�\���:G{:���9{�����ԍ�����d� �7{�`�P�&�.��`ԏ�o�o00%U6 �j	��o0�ۏT�?�x� c�������ү����� ��>�O��pO�u�$� ��9�����ڿſ��� "���X�C�|�gϠ� ���ϯ��������͟ ?������%߇��� ���������,��P� b�M��q��Y���}� �����:�%�^�I� [������������  ��$6!ZE~-� �Q�c�u�s�o  D/hS��� ����
/��./@/ ���v/a/�/�/�/�/ �/�/�/??<?'?`? r?]?�?�?�?�?�?\J�FEATURE �U�U�P	a�Handlin�gTool 'E �allyEn�glish Di�ctionary�-A, PaM�ulti Lan�guage (G�RMN) t\i�r4D St�@ard'F  p�rodAnalog I/OzG�  VLOA�Ag�le Shift�zHl.pc�@ut�o Softwa�re Update  \pk4�C�matic Ba�ckup+Cirp�k�Aground Edit @�-A�@uCam�era�@F�I�@D�PnrRndIm��C)E�@Pomm�on calib� UI S �@�@C�onQSPMoni�tor,B�@�@kPt�r%@Reliab��@,Bduct�Data Acq�uisoS,BAD �p�Piagnosx�A�A*D
PCV�P�ocument �Viewe{R.@w�c.�Qual C�heck Saf�ety[Q �Pl@E�nhanced �Us�PFrP.@E�NDI5@xt. oDIO kPfi�Tu *`F-bend`ErrzPL�RdTKf�gs  ckTo�Icr�@3` BWD�*DINT F�CTN Menu�`v�S�AM@�`TPw In�`fac�e~{`t\jG P�p Mask Ecxc`_@�EHT�`�Proxy Sv��T�A�QHigh-wSpe`Ski;T�dPcs@�P7`mm�unic�@ons4.@�P\)qur�`�`��I.P�`�A�bcon�nect 2EWIwncr�`str�P��VcsgeK�AREL Cmd�.XG�e�sRun-�Ti$`Env�WK^�`el +�@s�@�S/W-A�PLicense�S��Vetw�PZ`Bo�ok(Syste{m)*D   Q@�ACROs,r/�Offse�@HTMaH7`�@J��@ngQ@echStop�a�tpp�RPsiQ@i�Ub�K p.f�@MCix`�@�@'Gt`�Q@od�@witc=hzH93 R��pR��Q.E� R808�͆OptmڈPJ�͆�`fil�Vt �I,`τ�@gOw 03\t�PSB-T�`
S�IPCM fun�w�cF OY�v�pR/Regi�r=p�q�GaPri�PF`� �ELSE���@Nu�m Sell�  �oadx���"` Adju-p*DN@l@˕��J \j76�t�atu��Xx˕�Y � F`�`RDM R�obot>@sco�veGA im�R�emj�7anqG !|b?�Servo7`���,B!��SN�PX b�rzH59y6�`�CLibrFCN۔H55��@ {�P��〙`��o�pt�`�ssagI� �aTCP �C8�}K6��/I�m 1�p���MILIB!�.vyrLP�`Firm�B�'Gj7á�`�bAc�cP	U
��Q�TX�J��55�Telyn8�"�55 (���$A4�h�I)�`To�rqu�@imulyayQQ tph�@7Tou��Pa�q'G�P�� P�Qփ&�`e�v.  i�U�SB port �SPiPN`a�P P�
!1�nexc�ep��Y�n�S 9� R�i'G "L�`VCWQr8r/rp�ڰ"���P��\����@�ı��T��SP C7SUI��hc�P���XC��MA,`We�b Pl�.�ER �`�y�O{�p̀/��`0d�Qz`R�?�<ZyC�@e�GridD�play BAe��X�D�QJ�iR��.qJx���ԍ�AAVM��eIO`pNa�PAxy`�,B77����-ATX�PL�+CHCSB�9�-2000iB�/210 V b\>��Ascii�aΒ�LŐ�P��L�c�Up�lŐ'G���A���`opPBA 0���A�qhW�����1�`CE�`{rkJ�g R7P�PRUT����LQRT/KeybowA�Man^@v�:��PC�Pl sd�by 3E-c�Uol:@qQ#GuwF|�C�P�@�@�b�QkPss@tN@t^�� td\$�o�p�rE�s@�f ��LQyqc�@�r��ori`���P�PCS Jo��sc`����@��aL�Blu 4e��PH���<ZF�,`D�@in �N#ay�.�5LPDqy���ifi�SO 10i�`fDG@�p/�cUb�Outpu�B0�ࠃ`���oimiz��tm���KfAxis7a�Q ������fm��s�� w MS��FRL��am� ��P@HM�I Dev�p (��� ␠P�aΐ��{PM�h772��p.qnn/C֐o�ޑ�@J��x�oƃ #1��u��77�3.=��dЃZqRD��O���Qb����C�o�qTXY�RO�FINET�J "AM0�d�Dp��GRAM/JOG� OJ����@ ! ~d�Passwol�2i�R�`5!th�����8�SN�`Cli��Q#XM ��SPEE?D OUTP����c`�� RHi��s�=e801DpVAG�n�r��2"�!`vo�gi 7��BL$�#��3^.WeavI�~*���V��64MB �D <Z� Ġk2FR�Os;802DpAr�cҐviszS�*A�uxx�J&Celld�L6�9��OTsh�1(FM�@�<c݅]s�5��@p�  m�7t1y�@��@r2�@����(9���� � p�1`۔I���w�./s0��PR�� 2P���Q7� e�@`�LR�ZvE% �Pu+DDf(?�x��Pq`@5 f�T1G�T8���w 40� ���D�s��p,���t�BOPT��H�pQ�SN`�`cu��[Re� �p�S�yn.(RSS)z$QlU�quiry`�		 0��?����� �@8�t�
�QestbSm0t-ESS�L) ՠteHPWyS7@f��miLjECSp�a<_�N�h681�$r6'�dib� LJ���P cR��q��p�| iA/l��a71{a�p��=��!{aZ� �END  ��dpn����fd -�#V8.x I�(��!wEMZ$�EQ ñ�����LFRE+U �e��d@a1 �#�s\0� + ��� 8�when arg j�!����͡CD�tip*P=�Qk�͡u8sd �R.Skif�WF�,� BCK TseAb�v!a�ung�p�Ϡo�!r��PZ�!1�q68��I�Q��A F�`b.Ti�g/Td�(C� iox up�� l�b�of GOسT'o f��G�pQ�=m�psfmn�p��s�tQ� �:�-P+S-s�r�pL�@�A�ff.a.d S.�PN:FW-CHK JG"�� ���\cdcCD}:��SSTEP̢�BWD <�.E�r.af� 8x�Vag_C.l�j� ��tseJ�� Isms8` iq�+P�.Alloc.M�em.쀛k�29�P��� I����w .�K[�l Var.�Scr &�O|����FB_CMB�wlar��MNS�܏�I�wr.�!FU/NC-Mx�R9`���	s � S�˓k·n.sMP 6��Z��cmd.er..-Pdl.�Prp�8�aEC#rignǱ�&� f� }�TSHE�LL Hebe�at���No�.�On/��w.SRVO ?!���,�9�]m�� aw��6���GunM.DO.�@!.Gen.�A �R71l���?�.s�crn free�ze qP3�81+Inv9`i�g.��ch�pel�dpŁx ABC�&"g�p~�X '!.d���.uP�p.��a�r gex.�4�.��.abd ?PGPX  R`�:k�.��spddѐd4����p�� P}�<��۳3wp0տ��"F�r��Rd�/�rE�C)��sg.E��;�!aσ� Anyl}ϟ�R788���ä0W��������anlg����`\H	�+ӲPp%�G�IS� A�c�Ur^��
Y�yߞ��8 J6�߷�(Lin��S������o\aw�����ӿ�C��Pk=��eco<Y�{�wmleu���MH Dϳ�48 �H���MH����Txِ���d "F�#�\mht�3�b��:�[�"AP�w�h�tot���B����E3TU����ol$�.�p�����l Ef=�5o�csQ0�)�;���
4�'545`�:�Ip��x���H574`��J�2���fa����`��j� ��cenl������sH50��INT/ ��`-/�ķ�I/k#a�f/�z�55��-�Ĺ/�#9��/'52��/�0K��J?"MN�/�50��4�rH~?�2Z�!�?��u�4J6_P�?�2��?"t42�+D&0M%O;��pBO� "@O��a�zO�Bic���O�#0D�/81�O�CpJ�O�_']��"_�Ӷ�8�ENY_lo�rϼ?H-�_�1�O��R/��*�o#bx�Po��s! ���- VUo»�Roo8�ϯd2 J�o��Vi���A0d�o�Ds_�.f �f�ib���CLo/�_2�O��Mp�;?��}vm\cv���Yt�T�T��Egnai��?]�����O�taX_N_4/�a���a.@���cb_-������e��;�a�a���bsi@��w��ޡ ���dӟ1Vig|?�l/~/��r+�=���a�S�𯗟y
n'�9�F���|�G�nP��gί�ѿc  ѐͿ�� A��531l~wO�O3 R=ϫ�RS?��3 F�6E09 ��W��o�_P��dm@To¿H�Z�X/u� �� ��U�0����A���/x��_�SEND���3 RX�r6��ef3J9�Ϣ�AC4��8P�_��mnm�~0��.�x���CRL�*�'\sf�v61���Aj�/�6Y@i���fK��	�j<��ߌ����ND���1p�f��fe�(F�?k�)�e�DB/t�f���ZOƄW "H�O10�F��fe"L��5,9 �o�t\ha�����}���3Ttr��^�h6h�J�.z��ʕ
I%/���nd�hm��buDE��L?��F ���V6���4G.$`j_��rl���/��0u?;��/�?YSC(? :?#Ff��_�e��9O+�H?�u74TO�D7 ( ?�����	�O^�fL  feIn\/��gJ5_�onO�VJ351�O*VI)�_�D�sfm�_/E�_��e�8�~_xO48�O"a�d$��I@/&�mn��o�c� 4Z! j��o#sioF_X_5�9�?3t8.o ingI7�^p�o�t��$|��5P���!Lo�w (B�8O����PE�������}��o �Oȗ����l_�/"/<��a� nit�/�E�pl4_��!
�o�n|�Ƈ��e GL�JETX�:K����674=��߱N 9#`�n�gcr��/�0�~u�ɯ{d.p����3da���74�ﾯ�`�r�HG�q��2.@p�vu����/��\��~�  :��2��c.p�21�k��3"�ݱRS78"�= P�0�?J614��(��ATUP  �ONY�545��Y�6��s'�VCAM/�C�RI��=�CUIḞ�Y�28O���NRE� t.vA���_ ��`A�SCHO@���DOCVO� -^��DCSU� p���J60^��0��EI�OCw�NT��54�"�i�2��9�� S;ki�SETw�q���1�J7��921�@�MASK  K�207PRX�Y�s��7�9�O#CO{p�@1�3���8�áQ{pkmaY�Q��m�39�s���kcklLCHN�~=�OPLG�A.�J50~�r@I��HCR�PE�I�CS�j��`l��Ђ�KAR���J55^�rt FI�DSWo3�q�����q�f`nI�PR r����f����R��aU�CM���ӡP^�jЀT���f�9�1�v��L�1�f�����v�209���PRS*�́Y�9J�V�FRD����|��RMCN���93xR�n�|�SNBA�@w1\k��HLB��ME"��M���������q�2R�in'�TyCj�1�TMILC����A®�p= )�PA�б�A�TX�Pkrc)�EL��Y��Ү�tY!Y�8E�rcfX�0C�.��Y�95����95f�f.v|�UsECN���UFR����X�VCC��v \�wVCO��1.fL��VIP.�735.��SUIpL U���XФ�W#EBj��1�T��	к��2��g JT�C�G��sIGr��I]% PGS�3�% RC.�I�s��\�at��H89v�8��U1�X��@�H610.�Q�l�R7�]ӱRx��t�69���9����� "Cfp�61���J8��A0Fp��v��q�7R��j670�3^�"FSGY�8^��1��)6~���HA�4��΀�X�~�m�55v�f;tp$ J56����&��R5��7%��R7��tun0�9�8v���5e�U�82.��sgt<�5����/����0.�70\�$ R55~�979.��J76R�O�0���573��J96 ѱ���"��g��.�+T"0�6YF> ��4.�)p� J���p��9����� ��57 �5�A��~����\� ��^�b��]�� ���в�Iß���:V�5��tdf�����^���9ѵ�D06^�mch��"m�� ܂���SVMr�men��LIr���v��CMSF�V"� j�&��TY��6�IÇCTOj�U����s�gm��5����NN���K0f�mku8�O�RS���%8R�$8v��lwEXT6 r��F��I#OPI6 at� ����/�R6!!|� ��PRQ  ���8L���Sd2�w8�2f�I�ETS6 U�wSLM*�svg�!6i��52^��� �޾�iase)�OA2� �)�RAN�&��3��VA����IP�N6H@.�=�EZE8�0�  UPD~�%�fU�MC~�1�P1I��3E0}�3�@"�� �@~���@^���@�&��@����X�P1�
��B.�9� �Bf���T2"�I#�@��al`'��@����P2Q  �B��n�`�7P.���6R~�tol��P92}��P22v�#P2��m�sP&7P~Їkse��sP�?�P24^�Fpl�7P^���أP����S3U�kks��P27v�� ����P���B���P3l���P4�1hk��3P5}�P5iQsP5I�a�P33��gkdf=e���������3J���U���s'gkt=e2 D=e�����
=eI����k =e1"��������� �����>��f5B��AB Ve��e��e>���qB �e~A��1����2���2 ����e��e���� >eV!�e�A���B�����eJ!��tQ�f� �e�2Q��=R�uJQ��hst.Ev�v ��m��e�!��ft�P�v�g@�R����������n�����4$��  p=e"Z�<fak9�v|5�o orcm=e�"CC�U�܇cc �f���d9��f������@�e]��g/`�:hm�� �hlo����9�k
�T� ֟�}y����!0	�yfk�weyoY��ve�0���}���un<f�z����fsub��c�fccce�+��fE�W�i�{�v��������Ğv����뛍iY��
!s����� Di������f R�vT� "(�58��v� ��vcs/ "�:�� {ag˗925"����f26' �fr��E^j�4ᨖ "sDG�/�adg8v��on ��,vM��߄vr��q�?dse���:�di�����!\�e�d -=ee	��yf���fN-��f82 vs�I�[�m�8vāϷel�Ϯ���slb8vG��T���ST��/�l�0�B��f�L����p�dtHf����dg��b�����'��������dju8v{41h�g�w��4�f51�vi2����n��ro�f�stK�nat�f0���  �=e�3����PG`onwSpox�, P�8�n�OFT|�bp�feqi�f�v�alu�f"WE��<͌8vsweq���E�7`tpȦu "�p�&V�n�wvKq"�v��onf�v�z��ui��APF�@�΀�s��ftp �f����T������bw8vI�����&f��-\��OT�#/5-dvG/Y/k'Kc93P�/�k9P�/�/ "K���/��  H5�5
P�!I1!IK9C46!I�!I=a!I �1!I�Q!I�3!IA!I9!!I�05!Iq�!I i!�J�0!I9a!I�0PJp�!IaqJ"SC!IY11J�!IP� !Iua �J�!I�qZ�!I��8�Z�!Iin.@J�_we�_�_%V��1_X�p�_�Yu�J]_o[=o?[ld_o�[_Ko�_�_#Ghomj)�!Ig\ff!IU�1O#Gx��O#Gaxtd�O��O�o�oa��o�Yax �o'��4ASy�swas���#��ztp�J}1Q�h��FGMQOcG� �J-^h5 ZAR"8�k�0!Inrg�j-M�510�O_ė " �-�0\s`zyaJ���JMNI��Hf�mn��)1Z]���N�JP"q�cGmnm��Z�M^�0�~_�[t ���1���qOÏEW�T0Z�m�������P9D �]Mpsy����2dFFί�Zrl��0��0�FRA��`z�m��* E����er��ZM�_�RSo�1�y ������Ɵc� ��?K��CLPZ�}t�psZ]�o�PMA���Ims�J����n���ym���#�5�7��Y�낀�}��GRD0��]B��bd!�-R"�]�"�DN0!��"�odt`�-B"�-�"�=�r�P"�r^�"�-��"���"���"����S ��"��r"�n�i1�C��EM_�!�emd�������������� �
ssp
t� I)q"�asd�e!� !  � u�s@
rsal!�!w
IAR831din$�m�� Par��b�\�srg�F  !ޡ
! s�Se{rv�IF O��37 R�Loa�d�rvo�I)�o�R�def.z�s+! mi*GG C���0*8- x!+�Тng M�OE, P���A��gco��pL�migp*~F�*� �p�q�=0�f.s*h-��0e�NDO;�fd�+ -�+ivqe��²)691!:wRIN�701�pti*��2I�} �+j`:j703��* OpJ�?O!K3�set,!?�O�?d��+M� �:dnp*�ER J�1 R�6ZT_+ (MIn�voi@* "�+���?$H6�*g.f�@*Jog�R592��che@*^ � j�r�_Wog�*l�ink�k I/\Q_#H J5A;P0*w J8�j/O,�읂B)cl�*v
x�J~`�*pprx�J�ro0z�o�k J68o��B(�P :]��r/�(mPj��Si�mp�te�+R609�[L�z��o�Z�toPjspa*tc�h�Jth *AST� kHST�*794�zin�T��a?S{ta *��Aϋ���b��_�5pm.pJCP�|58�J�ModbAOSO�bt�;��+PROp [ �O"�930�;�/:30\0�_�+�FSW�}�o�h9�pZam����*t\�j�p J�? ��C1o/�]]=-ol/�N���=8\gpJ�0��&�RCo��e�Np4�}_i0*VM���_�[�0 j92o��P��ceN�:�M~P0:(�N?+ WC�O�)dnw�EN�:��w- L�I/F ksJ5��r w�:ar��rj?��}@�cm�n a0�M=.�0����U�g�r)�c�p* j6�TorP_R�D)��=o�OkM�CR HA� H�j�=1\�;�=�@8�*^�@*h f�z-�@��82 (a*r :���������\��P:982�*0�(0�B��'0_�Sq������������0��P:5�80�*1�\ paN��j����5�����We�mOkm�4��\n�-A���804� j΀ �usO�-�\0�ڍ�a*n p:�M,���ZJ9ϫiM !
@mq�M`q�p�zj~,moo� �����@��i7�J�� zm�/hcυ( l6�
H5;g806 �M�54_�9nN�`�cz\P����  ST�D��LANGK0-�1Em�C%E��%E�671%Em�%E w(SemFCha%EQt��%E�� %Ej]@P%EM�%E��6IG!�FC- wO)A-%ECmp�%EJ�HM�%Eg S�V%Eo H�F>�P"IGPHF�!%Eh�p�H��F���Fn�mFfunLIO�83`OrCt%Ectio�F=0%Em�%E83\s%Eq�G�83�H8�FD j%EutpumF] �G19UF9/@"U=�%E(`!V%`mF��%E�@pf846\%Em�mF�j84%Gg M90%EHiOpg2hm!x%E�%E00iA%Ept,�F�%E͑%Em94l%E��f>�p�fZ_l_~XInt�FNQI758�_
�FXf�rfaPV�_'C58�\Tv�k75�o��F�L-�O;�-��o�k-�ne�V=1RB�T
r�P_�9\f�0p_��S_��p9�OPTN�B5��S�afe��by F8��QB��586<@��6q��=љ����э��]��������!���r4��]r��ir��}R�� Tri�����o25 H��PRA�$���o�Q��r6Q~�C��NQ��gRq��]!���q����O��!A�� ��F�Q��j62ޘ�! ma��- �P��napȆ��96�iBZ�(;����\/�%�DPN)@ ��൥I���U���Plu�����B��7҂��݃ۤa��1����������pΒ���Ҭ�P��IZ�]���������R�754�k�I�0�bskl�����]�萷�i1^���sr�ts/A·�D]�妕���J9�1���!ƺ�CUS8a���g�itpl�g�p�g���g�sdm�g�Sys<@gþ���R SMe�J73�7��Qf�P��Ds�K�g���Ie���e�\�sy(���s���m�enueŎ���Da9t0�g�etw��Ŏ��740��i�g� �(DT�.bO���Pare�9rf�Er��Β g�=�g�I�s�n�s�� Upe�m�g�07\{���R72m�9ǁ^g�4 R8��7�p�R"m�E�7 (A$E�j�,E�>0
E�f�dE�in\P��RR�ascbE��BR-7 TOE�rts�%�zR�RD�R617E�01��j�R6��6�09��1�j�TQS]�fo`R�BR�B6��qs4���U�! c=nE�ContE�p�rE�m�R56 JxE啲RJ756E�lNO�Rc5PE�q���"q��nsvE�Ep� 5�� E�bdr th��iv��ْ���55���0����582��J���88��"OB��bO穒�淐�^�NQB$mb����v��B$h848E�2�a�� 48s�UbB&���9 E�H6�12E�w� (��250F]Y�j�f�
\s���N��i�wh61��200��N�R H����L�3��B/1ybB$��b�\]�b��ae:�GK� I/��E	�79�P�$iBj�(E�G]e��/$*gd�\gY�#�gd�cmy� C�'Tr�p 22�煒�4����4yclX&ack8�/?5t8&�$��0��U��er|��t��4�H��CVT��;KL�� PH(����L���`90�30��8>�^94ǀ^M�����:E3 � w ]$CL\�����9��$�]Zq@] 9M�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿�޿��99G�����$FEAT�_DEMO U�@�A�;�   �N�D�Vσ� zόϹϰ��������� ��I�@�R��v߈� �߬߾��������� E�<�N�{�r���� ��������
��A�8� J�w�n����������� ����=4Fs j|������ 90Bofx �������/ 5/,/>/k/b/t/�/�/ �/�/�/�/�/?1?(? :?g?^?p?�?�?�?�? �?�?�? O-O$O6OcO ZOlO�O�O�O�O�O�O �O�O)_ _2___V_h_ �_�_�_�_�_�_�_�_ %oo.o[oRodo�o�o �o�o�o�o�o�o! *WN`���� ������&�S� J�\�����������ȏ ����"�O�F�X� ��|�������ğޟ� ���K�B�T���x� ��������گ��� �G�>�P�}�t����� ����ֿ����C� :�L�y�pςϯϦϸ� ����	� ��?�6�H� u�l�~߫ߢߴ����� ����;�2�D�q�h� z����������� 
�7�.�@�m�d�v��� ������������3 *<i`r��� ����/&8 e\n����� ���+/"/4/a/X/ j/�/�/�/�/�/�/�/ �/'??0?]?T?f?�? �?�?�?�?�?�?�?#O O,OYOPObO�O�O�O �O�O�O�O�O__(_ U_L_^_�_�_�_�_�_ �_�_�_oo$oQoHo Zo�o~o�o�o�o�o�o �o MDV� z������� 
��I�@�R��v��� ����ُЏ���� E�<�N�{�r������� ՟̟ޟ���A�8� J�w�n�������ѯȯ گ����=�4�F�s� j�|�����ͿĿֿ� ���9�0�B�o�f�x� �Ϝ������������ 5�,�>�k�b�tߎߘ� �߼��������1�(� :�g�^�p������ ������ �-�$�6�c� Z�l������������� ����) 2_Vh �������� %.[Rd~� ������!// */W/N/`/z/�/�/�/ �/�/�/�/??&?S? J?\?v?�?�?�?�?�? �?�?OO"OOOFOXO rO|O�O�O�O�O�O�O ___K_B_T_n_x_ �_�_�_�_�_�_oo oGo>oPojoto�o�o �o�o�o�oC :Lfp���� ��	� ��?�6�H� b�l�������ϏƏ؏ ����;�2�D�^�h� ������˟ԟ��� 
�7�.�@�Z�d����� ��ǯ��Я�����3� *�<�V�`�������ÿ ��̿����/�&�8� R�\ωπϒϿ϶��� ������+�"�4�N�X� ��|ߎ߻߲������� ��'��0�J�T��x� ������������#� �,�F�P�}�t����� ����������( BLyp���� ���$>H ul~����� �// /:/D/q/h/ z/�/�/�/�/�/�/? 
??6?@?m?d?v?�? �?�?�?�?�?OO2M  )HHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t������� ��ο����(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ������0�   1�,�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&�
7�:�-�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO�&O8I�$FEAT�_DEMOIN [ :D�h@�3@}PDINDEX]K�lA�P@ILEC�OMP V�;���AkBKE��@SETUP2 �W�E�B��  N �A�C_A�P2BCK 1X��I  �)�MAKRO900�.TP:G_3@%�E_?Z&_c_:G�E1__UT1]_C_�_D�_y\2�_�_UT2�_�_1onoy\3ooUT3eoKo�o�oyU9H�lJ3@�@8u �(��^�� �)��M��q���� ��6�ˏZ�ď���%� ��6�[�������� D�ٟh������3� W��P������@�¯ �v����/�A�Яe� ������*���N��r� ܿϨ�=�̿N�s�� ��&ϻ���\��π�� '߶�K���o���hߥ� 4���X����ߎ�#�� G�Y���}����B� ��f������1��K�@�P�O 2�@*�.VR:���RP*�����#S����yUn�P�C��RQFR6:D��4��X��T|@ |�y�_@I�xV*.Fq�%Q	�<�`�STM ���" ��RPiPe�ndant Pa'nel��H�/��/�Pi/�
GIFs/�/��/F/X/�/�
JPG�/!?�?0�/�/q?��JS{?�?�RP73�?O?%
J�avaScript�?�/CS�?(O��O�? %Cas�cading S�tyle She�etsTO~P
AR�GNAME.DT�O�l�\�OUO�1��D�O�O	PANE3L1�O2_%�_[_��_2P_�_EW �_a_s_oZ3�_:o@EW(o�_�_�oZ4Xo��oEW�oio{o�D�SHELLp�A %+rCm���G�ZG_MENUE0-O�u�q��~�EEINGAB�J�%3�K�L������vSUMM_VA'G.D>?�O:���������yTPE_STAT:��;�S��y�����E;�INS.XM[ҏ�@���o��aCustom Toolbar ���yPASSWOR�D�oU�FRS:�\C�� %Pa�ssword C�onfig���G>�CONF1��]���Aǯ����,��yEX?TSERVOC�U��K�c�������UIO�_SET|��%��AϿ	���4ϣyVW?EMZROUS�e��S�kϑ��ϼ�K�AGV�UP[�m����ϙ� �@���d�߈ߚ�� ��M����߃���<� N���r���%���� [�����&���J��� n������3�����i� ����"��/X��| ��A�e� �0�Tf�� �=��s/�,/ >/�b/��/�/'/�/ K/�/�/�/?�/:?�/ G?p?�/�?#?�?�?Y? �?}?O$O�?HO�?lO ~OO�O1O�OUO�O�O �O _�OD_V_�Oz_	_ �_�_?_�_c_�_
o�_ .o�_Ro�__o�oo�o ;o�o�oqo�o*< �o`�o��%�I �m���8��\� n����!���ȏW���{��"��$FIL�E_D�� 1X������� ( �)
�SUMMARY.sDG#��MD:W����s�Diag� Summary�����
��SLOG@��p���۟�����sole lo��~��TPACCN��v�%^�����TP� Account�in=���FR6�:IPKDMP.ZI
�j�
� ������Excepti�on$�ի��MEMCHECK���������/�Memor?y Data����� �)��HADOW������)����Shadow� Changes�,�ߴ�O�)	F�TP���χϲ��1�mment T�BD��ܷ\+�)�ETHERNE�T��͎f���3ߪ��Ethernet� 3�figura�C�����DCSVR�F�ϊϜϵ߸�%�z� verif�y all��cĐ{e�u�DIFF��p�ߥ�:ﹰ%��diff<���f�z�CHGD11��*� Q�����9��}�2����C�� ��j���GD3p9� �2��� Y����}�UPDAT�ES. ��ЋFORS:\L7��Updates �ListL͛PS�RBWLD.CM�{ό7�N0�P�S_ROBOWE9L��g�:SMp�)��M��/Em�ail��aïcį���Տ����  /��$/�H/Z/�~/ /�/�/C/�/g/�/? �/2?�/V?�/c?�?? �???�?�?u?
O�?.O @O�?dO�?�O�O)O�O MO�OqO�O_�O<_�O `_r__�_%_�_�_[_ �__o&o�_Jo�_no �_{o�o3o�oWo�o�o �o"�oFX�o| ��A�e��� 0��T��x������ =�ҏ�s����,�>� ͏b�񏆟�����K� ��o�����:�ɟ^� p�����#���ʯY�� }�����H�ׯl��� ����1�ƿU������  ϯ�D�V��z�	Ϟ� -ϫ���c��χ��.� ��R���v߈�߬�;�������$FILE�_7 PRF �����������MDONLY� 1X�� 
 �q�H��l�� y��k���U������  ���D�V���z�	��� ��?���c�����. ��R��v��; ��q�*<� `����I� m//�8/�\/n/ ��/!/�/�/W/�/{/�?�/?F?��VIS�BCK#��2�*�.VDM?�?0F�R:\f0ION\�DATA\�?)2�0Vision� VD file �?�/OO3?AO+?eO �?vO�O*O�ONO�O�O �O_�O=_�O�Os__ �_�_d_�_\_�_�_o 'o�_Ko�_oo�oo�o 4o�oXojo�o�o#5 �oY�o}��B �f���1��U��������MR2_�GRP 1Y���C4  B�r�	 .�ҏ�πE�� E�@��������πOHcG�P&�L�u�S.�K�y
�?��J���π:G:��r�9{��~��Ag�  ����BH̃�C��NƕB��	�ҕ��΄���πo@UUU�UU���S�΁>t�>�S��=�h=����>�=���;b��B:�{eg:�sX:�+N:I9��2���V�����̃E�  F,D.�E(p�D�����0E��5�D�� =��<Əd�������� �����οϊ���:� ��_���nπϹϤ� �������%��5�[� F��jߣߎ���J�\� �߀�!��E�0�U�{� f��"���F������� ��A�,�e�P�u��� ������������+ (a�߂�d� ����'���� ������� ���#//G/2/k/ V/h/�/�/�/�/�/��_CFG Z��T �/5?G?Y?���NO ����F1747�36h?RM_CHKTYP  0��r���00��1O=M�0_MIN�0r�W���0��X���SSB3[��_ �
D�e; C)O8K��TP�_DEF_OW � m���PGIR�COM�0aO��UN�C_SETUP  ��%O�O�O�O���GENOVRD_DO�6}�mEU�THR�6 dUd�T_ENB�O ^PRAVC��\�7�0 ���_�/��_�_|O�_� �_(o�_Lo^o�_mo oo�oyo�o�o�o�o $�oHZ�o~�h�3ydQO�@1b���r��eB�8��^���
��;�.���N���^�F�C%���E�DYZor��t >0��x����B��͒�B���r�	�y���!�&���"�D�F�x���������k�ɏ珑����1 \�>��:�\�^����� ˯Ɵ����ܯ ��At�V�'�R�t�v����ѿ�ޯ����OG/RSMTkScrY�p��0w�m�x��$HO7STC21d�y�0'�Qa}U@k����1��k�172.26.�27.230���e��*�<�N�`�n�e��ϒߤ߶������� �e	cfg_fanuc���.�@�R� b��Eu���eB���� ���������(�s߀L�^�p�������9�	�anonymous������e�w� ���t������ ��=�(:L^ ���������� 9K]6/qZ/�~/ �/�/�/q/�/�/?  ?C/D?�h?z?�?�? �?�//1/3?Og/ @OROdOvO�O�/�O�O �O�O�OOQ?_<_N_ `_r_�?�?�?�?�__ )Ooo&o8oJo�Ono �o�o�o�o�__%_�o "4F�_�_�_� �o��_�����o �B�T�f�x�����o ��ҏ����Sew ���t��������Ο ��+���(�:�L�o� ��f�������ʯ?Ώ��ENT 1e����  P!a��  �	�F�5�j� -���Q���u������ �Ͽ0��T��x�;� ��_�q��ϕ��Ϲ�� ��>���t�7ߘ�[� ����ߣ�����:� ��^�!��E��i�� ��� ���$���H�� l�/�A���e����������QUICC0�����!172.�26.27.861G#���	�2�s��!R�OUTER��!�7`��PCJ�OG7!1�92.168.0�.10CAM�PRT�c5 x1���RT ���%/�NAME �!��!KJLT�VL211350�R01RS--K�U1�S_CFG� 1d�� ��Auto-started2�/FTP=��!T� V��/��??1?C?U? ��y?�?�?�?�/�?f? �?	OO-O?O��/�/ �/�O�?�/�O�O�O _ _�?6_H_Z_l_~_�O #_�_�_�_�_�_o�>o 	SM<��� �O�_to�O�o�o�o�o �o�_(:Loo��o�������� �2�D��ZC��o g�y�������Z�ӏ� ��	�,�-���Q�c�u� ����THC����'� I��4�F�X�j�5��� ����į֯��{��� 0�B�T�f���ß՟� �ҿ�����,�>� 	�b�tφϘϻ���O� ������(�s����� ���ϔ�߿��������  ���$�6�H�Z�l�� ���������5ߛ� Y�k�D���[����� ����������
. Q���dv�����4(_ERR f�F*��PDUSI�Z  \ ^w����>WRD �?�%:��  �backu�p�guest�Tfx��3&�SCDMNGRPw 2g�%� ��:�\ kD?K�� 	P01.o05 8�  �_�  � ��_]  Nw���� ���y����2; ����������|+-(�  ���v@<+/=&9����V���? ��S/�  
� � �s#� ��{/�j���(����S�#�� Uң/� 5n 9
S`��d/!/�/E/�2���1234567&�?��?�? �?O�?*OONO9O^O �OoO�O#;�O�O�O�O y?�?�?F_�OV_|_g_ �_�_�_�_�_�_o�_ 	oBo�Ofo%o�o__ )_;_�o{o�o, )bM�q����Io���(��_GWROU�h�	-0%�	�!1�cxz���B�QUPD?0d6��C���TYv ��� TTP_AUTH 1i�� <!iPendan�������!KAREL�:*$�-�?�KC�T�d�v�L�VISION SETM�ԟ��\J��ٟ� I�'��?�9���]�o�𼯓����CTRL� j���
 �#FFF�9E3ȯ8�FR�S:DEFAUL�T2�FANU�C Web Se/rver2�
�, >۬����Ŀֿ�����WR_CONF�IG k� �f2��IBGN_?CFG l���2\ @\ <#�-
~�BH|�C��?�4:�~�L�DEV��`��V�� IO� ma�I�EXD�AT n����E�XFLG���T�FIL o����O�TP pYݮaR!�B���R ���	�MERCATOR�!RECO�� "R�_ACHS��ISKTW*�V�,�V�� "SENSP���TXQ�99�0 	Kein7e 0�k h�\?%IBSC����,M�4�8�@�EW����T�LMTN�  ����  ���������l�X�OSBAD�� 7�^�xT�DL_�CPU_PCQ��\B�B��� A8;\�[�MINd�� =���T�GN���O�H���рIN�PT_SIM_D�O�����TPM�ODNTOL�� >��_PRTY�����Q�OLNK 1q�@9K]o����MASTE�����SLAVEG r���OZ��UOv �C�YCLu�$�K�_�ASG 1sY� ����a�՗�~Z���`�$0c� ������a������ �%/0/B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�NXNUM�����IPCH?��O_RTRY_CNQ��I�D�N؁��8�b� �Z�t�p�FO�T�SDT�ЧOLC�������$J23_DSP_ENB�0�ь@?OBPROC�C��n�	JOGI�1ukL��ad8�?P����O�??�ۯ4_�pQJ_o_�_�_R_ �_�_�_�_�zO�y8!�O-oo)_;_�_ �o�o�o�o�o�o&oJ�B1+oeN aoso�o������(�:�L�^�9���BA c��������� *�<���`�r�����q�����C����?�BPO�SF�OF�KANJ�I_� K���RE$_�.Av/��/���>��KCL_L��2��?�EYLOGG+IN7�М�����$LANGU�AGE �����ENGLISHY ١�LG-Bw �VS���S�x �����B����S�'� ����Z�MC�:\RSCH\0�0\Xﶠ��ISP x��؊�⍊�fߡOC���Dz����AݣOGBOOOK yYݟ$�챟Xx�	�� !�]�x���`͛ѧ��ه	ε��>���ϼ̲_BUFF7 1z(�ϟ��ߞ /��K�]� �߁ߓ��߷������� ��,�#�5�G�Y��}�������DCS }|ؽ =��͑� L���$�6�H�Z���_IO 1}cJO�������������� ����#3EWk {��������/Cn�ER_ITMhNd���� ����//,/>/ P/b/t/�/�/�/�/�/��/�/?��qSEVt@�mTYPhN��l?~?�?=��R�S�0����BFL 31~|�@��O�O(O:OLO^OpO�?T�P��y[2��NGNAM]��6ˢ��7UPSc�GI�0c�����A_LOA�DPROG %��%UP021�}O��MAXUALcRM�ܑ��筥9
DR�A_PR�Dܐ�³ڑDPCf��ع�ͪ_$�;Y�P_G�RP 2��[ ��S�2S�	[1�>ڐ+  ��_�� �R#oo oYoK�Go�o so�o�o�o�o�o�o *<`K�gy �������8� #�\�?�Q���}����� ڏ�Ϗ���4��)� j�U���y���ğ��� ӟ���B�-�f�Q� ����������ǯٯ ��>�)�b�t�W��� ���������ݿ�π:�L�/�p�[ϔ�=WD�_LDXDISA��@+;l�MEMO_{AP�@E ?�K
 T����߀�&�8�J�\�n�DPI_SC 1��M��� ���T�Q���߅���� 2��V�h���w�K�� ��������
������ R�d�O���o���-����������*��C_MSTR �,=~ISCD 1��������� �:%^I� m����� /� $//H/3/l/W/i/�/ �/�/�/�/�/?�/? D?/?h?S?�?w?�?�? �?�?�?
O�?.OORO =OvOaO�O�O�O�O�O �O�O__<_'_9_r_ ]_�_�_�_�_�_�_�_ o�_8o#o\oGo�oko��o:MKCFG ��X�ogLT�ARM_�b�X;�b �c��� (t�b_GRP_�DO �X�`�����L��uq>k������o$MMETsPU���b��`	�NDSP_CMN�T��`�Q  ��I��q�al�v��P/OSCF"��f���RPM!���STO�L 1�X 4=@�`<#�
���a �� �����"�d� F�X���|���П��ğ ����<��0�r�\���SING_CH�K  %�$MODAQ�c��o>�i���DEV 	>X
	MC:C���HSIZE�͚`����TASK %�X
%$123456789 M�_���TRIG 1���lX%�ܪ��c��Կ ����˿Ͽ�<���� 7τ�+Ϩϋ�aϣ���`�������/�YP����`��EM_I�NF 1�w� `)AT&FV0E0%����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ������H�����D���AL�t�/������� ����߸��� ��M� �q������Z� ��������%���� [� �2����h�� ����3�W> {�@�dv�� /�//f@/e/�/ D/�/�/�/�/��? ���a?s?&/�?�/ �?v?�/�?�?O�?9O KO�/oO"?4?F?X?�O |?�O�O6O#_�?G__�X_}_d_�_�nONIwTOR=�G ?���   	EX�EC1�c�R2�X3��X4�X5�Xp��V7*�X8�X9�c�RkB Od�ROd�ROdbOdb OdbOd%bOd1bOd=b�OdIbOc2Vh2bh2�nh2zh2�h2�h2��h2�h2�h2�h3�Vh3bh3�R��R_�GRP_SV 1݌q� (d�?I���I?2������n��?g"6+�Ze�B���~e������U7�_D@R����PL_NAME �!>�Y��!�Default �Personal�ity (fro�m FD) �TR�R2hq 1�����Y� ? 	 d��� ŏ׏�����1�C� U�g�y���������ӟ ���	��+�2��K� ]�o���������ɯۯ��<:��)�;�M� _�q���������˿ݿ��   ��\  �  ���  ��  A_�  B�T����
��
��@���  ����B��p��  C��C�P D�z  E;� E�@ D��c�C�J�q�X��d�Y�p� t�l�`�u�e���È�d�\�]�E/~ĉ�\�����`@o�e��`ż� �E	נŌ��^Ì��t�\�@�T�|���EZ��å�]�x|�Yũь� EY� �ߧө������¡���]����ө������� /�������� D�M�a���q�]����x���T�E� �� ����]��/���-� O�Y�M�s���������`������ V��4��D���ECvؕњ���r�(>P�d�tl~ c��! ����� ~q�� 'EKi����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?-�F?X?j?|? �?�?�?�?�?�?�?� O0OBOTOfOxO�O�O �O�O�O�O�M�� �O\)�_E_���c_ u_�_�_�_�_�_�_�_ oo)o;oMo_oqo�o R_�o�o�o�o�o %7I[m�� ���o���!�3� E�W�i�{�������Ï Տ�����/�9O� ]���k����!�� ����s!�C�9�g� ]�o����̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�??X�j�|ώϠϲ� ��������O�0�B� T�f�xߊߜ߮����� ����_�%_>�P�� t����������� ��(�:�L�^�p��� ��c��������  $6HZl~�� ������ 2 DVhz���� ���
//ן9�O/ ]����/���/�/ɟ۟ �/?��??'?9?W? ]?{?���/�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_?�X_j_|_�_�_�_ �_�_�_�_�S_0oBo Tofoxo�o�o�o�o�o �o�o��,7�P� t������� ��(�:�L�^�p��� ��c��ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟����� �2� D�V�h�z�������¯ ԯ���
���/9/K/ a�o/���/}����/3� �/ω?�?�?3�9�K��y�oϝϨ��$MR�R_GRP 1��������� � `� �o ������ @D�  ��?������?������@�T;g�Ũ���*�;��	l�	 �����X�'���F�O��^ �,X� �k���K���K��eK����K~o�K{GK�M�sA�S���߈��?�;g?�����@
����Р����I����
��}v=�����X����4  �p  ?�
=ô7����A��  >�L���������	�������Ѡ����(Ѵ��,  �p�  �2����������������	'� �� )�I� ��  ����:��ÈM�È=��9�e���@u�{� v���������������������@��?��@�t��@��@�)��C~6�B�  CfK �B�B��Q������CR��| �� ��� *�ވ� H�B<�� �� ����Dz��O��$�J!��� �qxy�jz  ȅ�:y�� ?��ffؿ��O G���,68��@/(*	ѝ�=$0(��V%P_(z��U�UԿ��>�33��6;���;aʤ;r��@;��;�?	�<$D���/��A��+���?���� ?fff�!?y&02A�5@�,%5iq1 �-��]?��|?�'A� ��?�?�?�?�?�?O�OAOSO>OwOhF5F� fO�ObO�ON?�O�r9�O+_�HD�� �E�J ��E9� E�04_m__j_�_ �_�_�_�_�_o�_o Eo0e��nm2o�o�O�o�XG-��G���G���*��8ŬNg�� B�'o $6<�*:��?���_s9�B�@����4��yA� A��t<� 	����7��[�F�����d�k�����1�Ķ<��k��C�����` Ca���j~���~�}�!� �5���CHf�CW��FB�1B-v��=���%������XR����u���z�����ę����A�P��Blz���X��}�sp��R��d�
Ák��BU(�������F<rѵ��JGp�@KÌH��? I%K�Ab!���L)-yL!�G�Kӕ#HP� �H�R����(��L&��J�3�$H㞀H���A��|�j�U��� y�����֯������� 0��T�?�x�c����� ��ҿ�������>� )�b�M�_Ϙσϼϧ� ��������:�%�^� I߂�mߦߑ��ߵ���  ���$��H�3�l�W� |����������� ��2��/�h�S���w��G�E*��~�C�?yټ���Ć�����CV��L7�\]G��t�_�(��`��,�%����1V���A3>�8!3A��vM_���v3�g��y�!�;�%D93ҵ������	/�-/,�C %P�"P_.na{o�/���/�/�/�/�+� �/�/(??8<�8?G?
n`8"�ta?#?�?�? �?�?�?�/mo'OOKO9K�QO[O�OO�K�O��O�O  �e 3��O�O__�9_'_]_kZ  2 7D��EVp�U��Z�B
��q
�C)��Aj@��_�jϜ�_lD� CD�0ov;j�_@�_zo�o�o�oj?`T�aZ��4jj��1jyVZ�
 �o,>Pbt ���������[��a ��I̿���Ld��2NA� @D<�U�?ϐ]� � `��a�j�A�XU�Ij��;��	la�\!��ો��e��0F��a������5���'��0Ci �P������_��?����ǟ��,nP�P���V_�z&'��9�G���k����+UUp�s�=��ͭ���Y�Ϡ�Rۯ�Z�&f���G�TY3�>��u0  '  [�e�Z�B�ס��E���@����R��ҿb�B�P<�� @�Q.�abCp!��Tϛ�x�cψ�χυ�j����  �j:v�a�`x#�a���
�߮� R�dۖ��0yߋ�>Ρ�P���������F�>Lס ���Ao ���4��e�QG�a��*�?fff?-�?&g��σ��Yb��]v� ]���[���L桄x�� ��5� �Y�D�}�h���p�������_ F�P ����7��X��* �&������ �-Q<u`� �����N/r ;/�_/q/�/�/4�/ �/V/�/�/?�/7?"?�R�_4�Qn�,?�? |=(�0�~?�?�?O�?  O9O$O]OHO�OlO�O �O�O�O�O�O�O#__ G_2_k_V_h_�_�_�_ �_�_�_o�_1oCo.o goRo�ovo�o�o�o�o �o	�o-Q<u `������� ��;�&�8�q�\��� ������ݏȏ���� 7�"�[�F��j����� ��ٟğ���!��E� 0�i�{�f�����ï�� �ү����A�,�e� P���t�����ѿ�ο���+�R7(�����M�_�I��mϣ� ���ϵ�������!�߀E�3�i�Wߍ�{ܶ5P%�P����4��� B����	�B�-�f�Q� ��u��������� ��,��P��߹��� �������������� B0Rxf����  2K�� *<N`r��������/p"/A�F/T*
 T/ N7�ߓ/�/�/�/�/�/ �/?#?5?G?Y?k?�Ҿt/��{J��4��� ���1 @D��  �1?��3 �� `?7 �27 A��X�5���? ;��	l�2��}��KC�0"K> F��a��?/.�?:&�uO �L> �8�ObO@/�O�O _�O%_]�0@J_XW0�x_��AЙ_�X8_�_U+UU�_�_=���okiS/`0�09oGh�R&f]oom�2�	�o6^u0  '�o�h�_�o_`x,�2ZO2�hB Px~ @�`�u�aEC���o��o������R�p&�4� K ��r:h&Nq~U��2�|j�|�� !�в�ċ�q8�pڏ�>.a�0�1�z2�$��L�">L7a��pA��=���;����s�2��3�2�p?fff?�p?&ǐ���t�2 �4�y�5��8=��� D؟q�\��������� ݯȯ����7���Ffp&�s�"���� ��2���뿆����3� �W�B�Tύ�xϱϜ� ��������~_,���S� ��t�ҿ��߿����� �ߔ�
���O�:�s��^���AfpA�����������ꈕ �o��?�*�c�N�`��� ������������) ;&_J�n�� ����%I 4mX����� ��/�3//0/i/ T/�/x/�/�/�/�/�/ ?�//??S?>?w?b? �?�?�?�?�?�?�?O O=O(OaOsO^O�O�O �O�O�O�O_�O _9_ $_]_H_�_l_�_�_�_ �_�_�_�_#ooGo2o koVoho�o�o�o�o�o �o�o1C.gR�vw(���� ��{�����'� �7�9�K���o������ɏ���ی�P��P�.��~O��xT� ~�i�����Ɵ���՟ ����D�/�h�S��� w���W���=���  �6�$�Z�H�~�l��� ����ؿƿ��� �.�  2��T�f�xϊπ�Ϯ���������� C�(�:�L�^�p߂ߡ��ߴ�
 �ߒ��� ����)�;�M�_�q����������o�{J������� @D� � �?�� � �`?��!��A��X��I� ;�	9l!��}�k�e�x%�����F���K������������� =�����=(aL �p�y���������z+�v+UU03=���m����&f�������u0  ' /'(K/vo/��.���/Z(B �/�.� @[ �%[!EC 0�_/?[/8?#?\?G?�EO0�?�7  ȒO2:�֮!�!�pW<�?�?n? 瀈O$KV18O0:OHJ> ��)�M:�?�O�/��c>L��V0A��O �?�O�?O3!��!�� ?fff?� ?&'PR?C_O4.�"Q.� M9�}_��_Va�8_ �_�_�_�_oo=o(o�aoso^o�oR]`F � �o�o�o�on_�Y �oK�ooZ�~� ������5� � Y�D����R���ԏ 2��n��1�C�U��O j�|������ӟ������A� A��� '�0��T�?��E�>� ����ï�������� �A�,�e�P������� �����ο��+�� (�a�Lυ�pϩϔ��� �������'��K�6� o�Zߓ�~ߐ��ߴ��� �����5� �Y�k�V� ��z����������� ��1��U�@�y�d��� ������������ ?*cN`��� ����);& _J�n���� �/�%//I/4/m/ X/�/�/�/�/�/�/�'=(y����?; 	???-?c?Q?�?u?�? �?�?�?�?O�?)OO(MO;Lv�P�BPN��{��/�O8�O�O�O _�O&__J_5_n_Y_ k_�_�_�_�_�_�_o �Oy�Co��LoNo`o�o �o�o�o�o�o�o�8&\J��w  2o������  �2�D�V�d���� ������Џ�o��
 ��]OS�e� w���������џ������+�{B4���{�J��$MSKCFMAP  -�� wv�D�E�  ]�ON�REL  qE�t��p]�EXCFENB��
r������FNCƯ��JOG_OVLIM��d�����d]�KEY��z��_PAN���-�)�]�RUN���]�SFSPD�TY�@Ȧ����SI�GN����T1MO�T���]�_CE_GRP 1�-�t�\��	��-� ?ϗOc��sϙ�PϽ� t϶��Ϫ��)��M� �q߃�jߧ�^߱��� ������7���[���P��H��l�]�QZ_EDIT��n����TCOM_CFG 1�j���)��;�
��_ARC_�âqE�UAP_�CPL_�դNOCHECK ?j� pE����� ������ 2DV�hz������N�O_WAIT_L�����װNUM_RSPACEg���=��7A�$ODRD�SP^�ѨOFFSET_CAR�����tDIS�rPEN_FILE��=���SPTIO�N_IO#�5��M_PRG %#�%$*/".�WO_RK ��ԣ� G@S%��mDNC� ��m ��m!	 ���m!<�����TRG_DS�BL  -����z��/��ORIEN�TTO����C�선s�A rUT__SIM_D�q��D�TVXLCT ��#B�@-5_P�EXE�g6RAT�s0	�ѥx�k2yUP� �<>%�.����?�?�?OI�$P�ARAM2೏���&3	 d��VOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_���_�_o #o5oGoYoko}o�o��<�_�o�o�o�o &8J\n��}��x�����  ���  ��  A��  B�p��B���3�pH�p��  ���p�pB��pp�p� 0�!(�P� Dz  E;�� E@ D���C� 0��q�� ��p��������)�+���r �E/�!�,��qc�p���@������_���E	��C�/���/���������q���EZ��n�H� ���uL��� E�qX�J�L�t���0;�D�p� ���n�L�c�p���� ғ���� p�d������d��� �(�:�L�L��qE� �������� ��� ҧL�Я��q��(� :�L�^�p��������� �o���p���3���!��D�R� ĽĽ���p�� �� �Ϧϸ��������.� DO]�o߁ߓߥ߷��� �������#�5�G�Y� k�}�������_�� ����1�C�U�g�y� �����o��������	 -?Qcu�� �#1�x��0��}� <�*<N`r �������/ /&/�J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?9/�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�Oi�˿ ݿ�O�_%�_M_[� �OϘ_�9���_�_ �_oo/oE�^opo�o �o�o�o�o�o�o  $6HZl~�� ������� �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������� ���?�*�<�N�`�r� ��������̯ޯ�� �&�8��\�n����� ����ȿڿ����"� 4�F�X�j�|�K��ϲ� ����������0�B� T�f�xߊߜ߮����O �O��_C_)�7_1�[_ m_�ߘ���-o����� ������Eo��p��� ������������  $6HZl~�� ����� 2 DVhz����� ���
//./@/R/ d/v/�/�/�����/۟ �/��?*?<?N?`?r? �?�?�?�?�?�?�?O O&O8O?\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_KO�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o{� ���C�)7�!_ m��o��-�?�)�������A��q�$�PARAM_GR�OUP 1��gX���L�`8� ߐ ��q~�� @D�  ��?�����?�p���q�C>�����t� � ;�	l��	 ����?�X�΀π����^ �,�X ���pH���H�ffH��  H��H�?WH-���|�#��o�oi���qB� ' B��������������s�4  �p  �
=É���������ȟ�sA�8�¼r��qO«�C���r,��2���G��wρ[��|�,  � � � ������M � Д�����u	�'� � Т�I� �  {��l�=��������@�"����F�������[�i�F����������CݐB���f������б���Ŀֿ�   ���CR>���� :��<�H�wB��L�+�Xŷ� 3�tŕqDz������Ϧ�����Ȯ��� �x ��!� � �,�:˅�!~D� ?�ff{xR�d��� ��������8�����ڰ�D�$����(����P�!��A�����f�>�33�}���;��;a�ʤ;r�@;���;�	�<c$D4�q��A�s�ʴ���?3�q�?f�ff��?&����A����@�, ����©ᵄ�ɤ�� ��#���脃�X�C�|� g��������������� 0T?x�����q�mD�� �E��j E9� E�0�&J 5nY�}��� ��{�-�:/�[/ ��/��/�/�/�/{���?��|�3��BA��/=?(?a?L?�?p9A+�A�4㠰1��?��y?�?u?O�<?��OOKO6OaIm���k^OC����` Ca[OH*%D�%@$A�A@I��ܾ��CHf��CW�FB�1�B-v�=����̞�����XR���u��!_DA�ę�����AP��Bl?z��X��$_0���R�d�
���k�BU(��无����E@K����JGp@KÌ�H�� I%K�A	�aLL)-y�L!�GKӕ#�HP� H�R���_�P(�L&���J�3$H��H���A��_ #_o�_5o oYoDo}o ho�o�o�o�o�o�o�o 
C.Syd� �����	��� ?�*�c�N���r����� ���̏���)��M� 8�q�\�n�����˟�� �ڟ���#�I�4�m� X���|�����ٯį֯0���3��G���b��%�C�?�c�j��������CV�a������޿��@��O�:�s�^�(d�g�`���0�����dų1V�Ϯ�^��3>��������v��߰�v�3�g� �2�!��;�%D93ҵ�L�Lٌ�z߰ߞ���\��^� Pl�P�!"//��;�e�P���t���������������8�0t ���S�>�w�b���B�`/�����������08&HO�HZ�  �e 3� t6����  2 D�7�E� 1���B��1�1�0C��@��A���@�?z���D� D��������/!/3/E/W/���?�p!����R������� ��
 ^/�/�/�/ �/	??-???Q?c?u?��?�?�?���! �����̿����tK�&��1 @D�0��1?vPA � `�V�By��4�1�2L;��	lB���RKLC@iK��F��a�2O�?�O����O��L��Ci�O�O����i&_��J_5_n_YZ,��@�_�V��_!��A��_�Xa_o]U�+UUoo=���Tofk cv`�0�o�hb&f�o�m�2�	�o>U^u0  '��v`B�~a)�oM@_H�B�OyAxBU<��| @e�t4C�F�B�
��C�.�,b6�m�{�  �6�:�"�!� ��B>���ÏU� �����=�+� �2�>ua�0V�=�y�k���I�>L~a�T=�A@�����ۏi%	A�3|B�p?fff?�p?&�9�*�6�B	� D4�Ed�H���HD �����ܯǯ ��$� �H�Z�E�~���g��� ��ؿO�q�s�ѿ2�Ϳ V�A�z�eϞωϛ��� ��������@�+��_ s�9ߚ��������U� ��*�<�۟Q�c���@���������T��Q_��8�#�ϕ �o%���q��������� ����(L7p �m������ �H3lW� {�����/� 2//V/A/z/e/w/�/ �/�/�/�/�/??@? R?=?v?a?�?�?�?�? �?�?�?OO<O'O`O KO�OoO�O�O�O�O�O _�O&__J_5_G_�_ k_�_�_�_�_�_�_o "ooFo1ojoUo�oyo �o�o�o�o�o�o0 T?x�u�����w(�q��� ���&��J�8�n� \�~�����ȏ���ڏ����4�"�]�P̒Pf���b�����x�� ş���ԟ���1�� U�@�R���v�����ӯ ������`�*���3�5� G�}�k�����ſ��� ׿����C�1�g�u�  2�ϭϿ��π������+�=�K� ��o߁ߓߥ߷��������
 ����D� :�L�^�p����������� ��b���o�{J�_�+��[�H� @D� � \�?�b� � #`?��h���C]�\�|X��� ;�	lh�c�}�����l�����F�������+����.�Є�N 	�߄o���� ]�����]�Y�.��@N�r�+�UUwz=��� ��`�X���a&f/-N�[�:/�?u0  '`/n( a�/��/�u��/�(B �/> 1@� 45�!ECw��/�[?�/?j?�?�?���0�?�7  Ȗ2:H�S��!%h��<8O#O�? .�YODkK�18�0�O�J>��I�p�:�?�O�/)�>1L�Sĝ0A��ODO�O<O�3h�N�h�10�?fff?40?& nP�?�_�4u�iQu��9 d��_b��_SV��_o o<o'o`oKo�ooo�o �o�o�o�o�o�o8 �_�_�_1�-�� �����4��X� C�|�g�����%ӏ�� ��U�yB���f�x� ����;_��ß]���៰��>�)�A0A�f��n�w�6����� /U7/���ѯ
���� @�+�d�O���s����� п�Ϳ��*��N� 9�r�]�oϨϓ��Ϸ� �������8�J�5�n� Yߒ�}߶ߡ������� ���4��X�C�|�g� ������������� 	�B�-�?�x�c����� ��������> )bM�q��� ���(L7 p�m����� �/�/H/3/l/W/ �/{/�/�/�/�/�/?��/2?7($1���T?f;P?�?t?�?�? �?�?�?�?�?(OOLO@:OpO^O�O�L��P,R	P�N Q¤%?�OI8 �O%__I_4_m_X_�_ |_�_�_�_�_�_o�_ 3ooWo�O���o䈓o �o�o�o�o�o% I7Ym����w  2Ro��� 1�C�U�g�y��������Ϗ����)�8HoM�[�
 [�9� �O������П���� �*�<�N�`�r��B{����{J����􋐻B�� @D��  ��?�£ �G `?>�Ȣ>�C������F� ;�	lȢ�A}���̠<)�E�F����6���A��|���E�� ��i�G��Ͽ��,� ͽ� �Q�_ǽϹv��РϮ�!�����+UU����=����&���6и�@�N���&fd�vݮ��y��~=�u0  '�� ���������բa��9��B W�� c@����EC�A ������������q��-�;�  ���:o��qU��uȢp��q���� �@�������8������> 5ѩ�С��9�+Sc>L>ѳt��A�D ��B����Ȣ��Ȣ���?fff?��?&� �����բ�դ ��ĥ$¨D��� xc������ ///>/P/'/t/_/ �/13�/�/�/? ?:?%?^?I?[?�?? �?�?�?�? O�?��3O �?ZO�/{O�/�OO�O �O�O�O�_#_�OV_`A_z_e_�_�_Am�A��T��S�_�_�_ �Z����_Fo1ojoUo go�o�o�o�o�o�o �o0B-fQ�u �������,� �P�;�t�_������� Ώ���ݏ��:�%� 7�p�[��������ܟ ǟ ����6�!�Z�E� ~�i�������دï�� � ��D�/�h�z�e� ����¿���ѿ
��� �@�+�d�Oψ�sϬ� �����������*�� N�9�r�]�oߨߓ��� ���������8�J�5��n�Y��}�(��������������
� ��.��>�@�R���v��������������eP�P&=A"d��V ��[�p���� �� K6o Z�~�^ O�DH ��/=/+/a/O/�/ s/�/�/�/�/�/?�/'?7  2�[?m? ?�?�?�?�?�?�?�?JJ?/OAOSOeOwOp�O��O�J
 �O �G�O__0_B_T_ f_x_�_�_�_�_�_"��O��{J��$�PARAM_ME�NU ?�U��  �DEFPULS�E�[	WAIT�TMOUT/kR�CVBo SH�ELL_WRK.�$CUR_STY�L-`nlOPT�A9a�oTB�o�bC�ioR_DECSN :`�l�o�o1, >Pyt�������	�aSSREL_ID  �E�1��USE_P�ROG %j%8�j��CCRF`*��1c}�_HOST7 !j!�����w�T7 ��ۃ�����݃�v�_TIME�Db*���`GDE�BUG(�k�GI�NP_FLMSKl@�o�TR~� q�WPGA�� _��I� ���CH}� { q�TYPEl@��4�]�X� j�|�������į�� ���5�0�B�T�}�x� ����ſ��ҿ��� �,�U�P�b�tϝϘ��ϼ���q�WORD� ?		FwOLG-c	U�	MAKRO+�_SUCHL�C2��S7T�TRACE�CTL 1��U�a
 0' �(�@ U V�{�2�ߗߩ�S�D/T Q��U��o��D � 	� �`�а`���` ��'���-`��F��\�*��H��I��J�����B���M���`��6Ј��7 ��Q�ԝ���S���F`��U��V��W���X��Y��Z��[���\��]��^��_���`��a��b��c���d��e��f����<  	� ]���� �#��#�U�#��#��#��#�5�#�����r���!�1m��Pm�k�z�(n��n�k�k�j�U	k�
k�k�k�k�c���g��g�^�� ?��@c�-�q��	����`�������
��	�9z�? ��? ��?  ��? ��? ��? j�? ������� ��_�	_I_Q_Y_�i_q_y_��_
��_��_�� *��U��c�l	UlIl���q��y���)��ؑ�ؙ�ت���i�ر�ع�ت�����������l*Ylali `d�Um	mImQmY�mam��1� �q��z�����P#������q��y��Ɂ��!&��ə�ɪ���i�ɱ�ɹ��*��������������������
��D���Ժ����U��������Q���@������Q��ސ��!��"��U#��$��%��&��U'��(��)��*��U+��,��-��.��U/��0��1��2��U3��4��5��6��U7��8��9��:��U;��<��=��>�� �������/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OL ������/�A�S�e� w����������� ����/�/�/9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�	//-/?/ Q/c/u/�/�o�o%C�e o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� �ek����� %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o��o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�����/�A�S� e�wωϛϭϿ����� �����o=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?1�?�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y�����s?��ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� ���������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o�� 1oWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c��u��$PGTRA�CELEN  �v�  ���A`ȋ�_UP �����������y����_C�FG ���T��Aa������Ā�����������D�EFSPD ����@a��Ћ�I�N��TRL ������8��V�PE__CONFI����ş������#�LID�á��~��GRP 1��� �v��CH������AaA�  G�G� G�7�F�,� A�  D	���A`d��)�9�~��� 	 �8���S� ´��n��B����������������B>Áe�G�Y�C� <,1<49X^� ��Z�����������v�� 9��IoZ�z�����
 B�������^�m���A��G�?��G{l�| �� %K6o�Z��>V�>V�z�v����/^�!��
V7.10beta1�� @�33@�2�\@;�C�RA`C C>  C�W��T#D�� �j"0�g!����� Dj\ 2 ��BY�\ S C] �p����!,�!p�A����Ak33>����B �!@�� ��ffA����@������ ���K�'y`T"���/?���&�8�ѩ��[?�? j?�?�?�?�?�?�?�? !OOEO0OiOTOyO�O �O�O�O�O�O_�O/_ _,_e_P_�_ܳ �_ �_n_�_�_�_oo=o (oaoLo�opo�o�o�o��o�o�./T#F�@ >y:}N`|~ ?�&������/ �??/?A?J��on� ��k�����ȏ���׏ ����F�1�j�U��� y�����֟�ӟ��� 0��T�?�x����_�� ��o��ϯ��,�� )�b�M���q�����ο ����1c=�O� y���ϸ������ 	��-�?�H��l�W� ��{ߍ��߱������ ��2��V�h�S��w� ������������.� �R�=�v�������[� ��������*N 9r�o���� ��/�a�;Mn��ϒ�����$P�LID_KNOW�_M  :%��>!�SV g���������)/;/ M/�q/\/n/�/��� �M_GRP s1��� lCR�"��� ��&�$ �0H��@�("1*5&?8< ���	7�+a????�? S?e?�?�?�?	O�?�?�9O�?OuO+D�MRJ�#��-T��C5��"�C�� ��O �N_�O���O>___ $_�_H_�_�_~_�_�_��%ST�!1 1���"`� 0�EZ�_������^�m��A���G���G{l����FvoYoko }o�o�o�o�o�o�o MCU�y����o2o)`� �C��8�J�x�n� ����ӏ��ȏڏ��� �"�c�F�X�j����������k3�(�� ̟-�n�Q�c������� ��������4��)� ;�M���q���Ŀ������c4�'��˿,� m�P�bϣφϘϪϼ� ������3��(�:�L� ��p߂��ߦ߸���c�5�&���<)�n6�%�7�I�cA7b�t���c8���������cMAD � �$"c  �dPARNUM  ��"�!��7�_T_SCHN� \��
��o�����UP�Do����S_C�MP_� Q���'��S_ER_C;HK6���cO3ERS�@��"G_MOP���_���RES_G`�z� ?aC�v�BS�SH���EI�r�OOUL 16gZ�~�� ���	/�-/�� �1//�/y/�/�/�/ �/�/?�/(??L??? Q?p?6/��Q/�?u? �?�?	O�?-O O2OcO VO�OzO�O�O�O�O�? ���?�O�OD_7_h_ [_�__�_�_�_�_�_ 
o�_o.o�O��\_Qo�a�no�o�o ���o�o�o����ox�V 1������ �^�`��^h�]�T�]���THR�_INR� S��dz�d�vMASS�� Z�wMN��sM�ON_QUEUEG �š��ȡ�u%MJ� 2��y���4A�  Y@�߉�Bʡ�!U	�N- UqN�v_m�ENDo�����EXE������BE���y�j�OPTIO�v��m�PROGR�AM %�z%�l�J3�k�TASK�_IP�ߎOCFG� ������OoDATA�1�}�@ 0��2 ޟ����&�0�ڑ ; &F� H�Z�l�~���B������������է�ׯ��5P�  ڟ*�<�N�`�4�����������Ͽ������)��?�G��� �j�|ώϠ�t�Կ��)��������;�9�0=�A���a�Gá�A� �Ϯ�������8��� ��5�G�'�+�]�u�Y�x��}�s�INFO���}���#
� �.�@�R�d�v����� ����������*�<N`r��I����� =is���DIT �}�@mU��>��WERFL��rs���RGADJ ��}�A�  '?���3�qm�x��~U�?C��@��<@�����%�qq���I�J���U˒��\9f�qrbbA<t�t]$&* /" **:""��/'#2UL"G%��!Q)Q���q/sE/W/ i/{/�/�/�/�/�//? �/??�?�?S?e?w? �?�?�?�?�?�?�?O O+OUOOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_�_�_�_�_�_ $o�_�_�_oko5oGo Yo�o�o�o�o�o �o �o�o;1CUg �������� 	��-�?�Q�c�u������ 	��,��P� ;�	)u�#A���=�Ɵ ���
//�@/ʏ ܏q� ���L�^�˯�� �������ܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� Dϱ�h�zόϞ���� ������N��.�@߭� d�v߈ߚ������� ����*�<�N�`�r� ������������ �&�8�J�\�n����� ��������G��" 4�Xj|���� 
C.l�v<� 8�؟���� �2� �����>/P/b/ t/�/�/�/�/�/;?�/ ??(?~?L?^?p?�? �?�?�?�?7O�? OO $ONOHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_o �_�_�_
owo.o@oRo do�o�o�o�o�o�o �os*<N`� �������� �&�8�J�\�n����� ���#��G�^h�� ��R���ş�� /*/ �6/��ҏg�����B� T�~�x���������ү �����,�>�P�b� t���������ο�M� ��(�:ϧ�^�pς� ���ϸ�����I� �� $�6ߣ�Z�l�~ߐߺ� ����������� �2� D�V�h�z������ ������
����@�R� d�v�����������& ���<N`r ���� 9Kb��l���.���$�PRGNS_PR�EF ��W�� � 
��IORITY  �ݔ�����MPDSPON  ݖ���#�UT&�5&ODU�CT_ID �"��OGG?RP_TGL$m&�V&TOENT 1��i*�(!AF�_INEE �/��!tcp�/��!ud�/�!Oicm!?�Z"�XY_CFG ݸ�+ ��)�a #��?�?� ��? �?�5�?�?�?!OOO WO>O{ObO�O�O�O�OH�O�O_*Y#t3��� %�O_a_�>�) ��#�/�:_į_��-%�X�A����,  ����_
oo.o)(T�����0"�PORT�_NUM#� �%�_CART�REP& {<�SK�STAE' �jS�AVE �i*	�2600H60%1��!�_'3?K 	ox����ݓe������
�|JU��e]_�  1��+ p �2݈���#�������a_C/ONFIw0�Zg#��]�U�ޔ��0��בVȃPt22� ֋���[��C�U��$��q�2�։�a���UQ8��?�?&M��?V?Q����N���&n�=���?����RC���C�xXD�M�T������ɹ�U���l���Ř�ѐ�YՕٖ|V)#�V�p�� 凭 ����y���i����� _������_��U]�� A���Q�w��ۯ���� �#����Y��=�˿ )�sυ�׿鿻���� ���U���9�Kߝϯ� �ߓ��Ϸ�������� ��c߭�G�Y��}�� �ߛ����)�s��� ��C�U���y�����k2�S_MOTI$ 2�֋
�?���_@��);M��`�5����x����Z+= Oas����� ��y��#�&/./ @/R/d/v/�/�/�/�/ �/�/�/:�/7?I? [?m??�?�?�?�?�? �?�?O
??EOWOiO {O�O�O�O�O�O�O�O __/_*O<Oe_w_�_ �_�_�_�_�_�_oo +o=o8_J_Jo�o�o�o �o�o�o�o'9 K]Xojo���� ����#�5�G�Y� k�fx���ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����������)� ;�M�_�q��������� ��Ư���%�7�I� [�m�ϑϣϵ����� Կ��!�3�E�W�i� {ߍߟ߱��������� ���/�A�S�e�w�� ������������ �=�O�a�s������� ���������"� "]o����� ���#50B k}������ �//1/C/>Pb �/�/�/�/�/�/�/	? ?-???Q?c?^/p/�? �?�?�?�?�?OO)O ;OMO_OqOl?~?�?�O �O�O�O__%_7_I_ [_m__�_�O�O�_�_ �_�_o!o3oEoWoio {o�o�o�o�Q�Q�Q�e��i%�f�o�fEL <�o  '��m�c<�S�e  8R�Q8_���� �_�_� 	��-�?�Q�c�u��� ������Ϗ�_��� )�;�M�_�q������� ��˟ݟ����%�7� I�[�m��������ǯ ٯ�����
�
�E�W� i�{�������ÿտ� �����*�S�e�w� �ϛϭϿ�������� �+�&�8�J�s߅ߗ� �߻���������'� 9�K�F�X߁���� ���������#�5�G� Y�T�f�x�������� ����1CUg yt�������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ ���/�/??%?7? I?[?m??�?�?�?�? �/�/�?O!O3OEOWO iO{O�O�O�O�O�O�? �?�O_/_A_S_e_w_ �_�_�_�_�_�_�_�O _+o=oOoaoso�o�o �o�o�o�o�o�_o "oK]o���� �����#�0 Y�k�}�������ŏ׏ �����1�,�>�P� y���������ӟ��� 	��-�?�Q�L�^��� ������ϯ���� )�;�M�_�q�l�~��� ��˿ݿ���%�7� I�[�m��z������� �������!�3�E�W� i�{ߍߟߪì����Ղ��%��������� ��%���Ӡ��� � (�B��8�O����� �Ϯ������� /�A�S�e�w������� ��������+= Oas����� �����'9K] o������� ���5/G/Y/k/}/ �/�/�/�/�/�/�/? //C?U?g?y?�?�? �?�?�?�?�?	OO? (?:?cOuO�O�O�O�O �O�O�O__)_;_6O HOq_�_�_�_�_�_�_ �_oo%o7oIoD_V_ h_�o�o�o�o�o�o�o !3EWidovo �������� /�A�S�e�w����� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o�����������ğ� ���#�5�G�Y�k�}� ������ſ��үҿ� �1�C�U�g�yϋϝ� �����������-� ?�Q�c�u߇ߙ߽߫� �������� ��;�M� _�q��������� ����� �I�[�m� ��������������� !�.�@�i{� ������ /A<Nw��� ����//+/=/ O/a/\n�/�/�/�/ �/�/??'?9?K?]? o?j/|/�?�?�?�?�? �?O#O5OGOYOkO}O@�O�3�1�1�E�I%�F�O�F���O�O�Ox�E�3�E  _2_�18?_u_�_>�_� �?�? �_�_�_oo1oCoUo goyo�o�o�o�?�_�o �o	-?Qcu ������o�o� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ�����
�3�E� W�i�{�������ïկ ������*�S�e� w���������ѿ��� ��+�&�8�a�sυ� �ϩϻ��������� '�9�4�F�Xρߓߥ� �����������#�5� G�Y�T�fߏ����� ��������1�C�U� g�y�t��������� ��	-?Qcu ��������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ ���/�/?!?3?E? W?i?{?�?�?�?�?�? �/�/OO/OAOSOeO wO�O�O�O�O�O�O�? �?O+_=_O_a_s_�_ �_�_�_�_�_�_o�O _9oKo]ooo�o�o�o �o�o�o�o�ooo 0oYk}���� �����1�,> g�y���������ӏ� ��	��-�?�Q�L�^� ��������ϟ��� �)�;�M�_�Z�l��� ����˯ݯ���%� 7�I�[�m������������%����ʹ��� ~h���������  �"ς�8�/�e�wω�� |��������� ���!�3�E�W�i�{� �ߟ�r���������� �/�A�S�e�w��� ����������+� =�O�a�s��������� ��������'9K ]o������ �����#5GYk }������� �C/U/g/y/�/ �/�/�/�/�/�/	?? /(/Q?c?u?�?�?�? �?�?�?�?OO)O$? 6?H?qO�O�O�O�O�O �O�O__%_7_I_DO VO_�_�_�_�_�_�_ �_o!o3oEoWoiod_ v_�o�o�o�o�o�o /ASewro�o �������+� =�O�a�s������� ͏ߏ���'�9�K� ]�o������������� ����#�5�G�Y�k� }�������ů��ҟ�� ��1�C�U�g�y��� ������ӿί��� -�?�Q�c�uχϙϫ� ��������� �)�;� M�_�q߃ߕߧ߹��� �������� �I�[� m����������� ���!��.�W�i�{� �������������� /A<�N�w�� �����+ =OJ\���� ���//'/9/K/�]/o/z|r�%�)%8�&�/�&�/�/�/�%p�%  8�/?r8?U?|g?y?� l ~�?�?�?�?�?O#O 5OGOYOkO}O�Ob�? �O�O�O�O__1_C_ U_g_y_�_�_�_�O�O �_�_	oo-o?oQoco uo�o�o�o�o�_�_�o );M_q� ������o�o� %�7�I�[�m������ ��Ǐُ���
�3� E�W�i�{�������ß ՟������A�S� e�w���������ѯ� �����&�8�a�s� ��������Ϳ߿�� �'�9�4�F�oρϓ� �Ϸ����������#� 5�G�Y�T�fϏߡ߳� ����������1�C� U�g�b�tߝ������ ����	��-�?�Q�c� u������������� );M_q� �������� %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ ���??/?A?S? e?w?�?�?�?�?�?�? �/�/O+O=OOOaOsO �O�O�O�O�O�O�O�? �?O9_K_]_o_�_�_ �_�_�_�_�_�_o_ _GoYoko}o�o�o�o �o�o�o�o1,o >ogy����� ��	��-�?�:L u���������Ϗ�� ��)�;�M�_�j�l��b�x���%s�����N� ]��͟ �{�����`���  8��b�8�E�|W�i�� \� n�����˯ݯ��� %�7�I�[�m��R��� ��ǿٿ����!�3� E�W�i�{ύϟϚ��� ��������/�A�S� e�w߉ߛ߭ߨϺϺ� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ��������������# 5GYk}��� ������1C Ugy����� ��	/(Q/c/ u/�/�/�/�/�/�/�/ ??)?$/6/_?q?�? �?�?�?�?�?�?OO %O7OIOD?V?O�O�O �O�O�O�O�O_!_3_ E_W_ROdO�_�_�_�_ �_�_�_oo/oAoSo eowor_�_�o�o�o�o �o+=Oas ��o�o����� �'�9�K�]�o����� ����ۏ����#� 5�G�Y�k�}������� ����ҏ����1�C� U�g�y���������ӯ Ο��	��-�?�Q�c� u���������Ͽ�ܯ � �)�;�M�_�qσ� �ϧϹ���������� �7�I�[�m�ߑߣ� �����������!�� .�W�i�{������ ��������/�*�<� e�w������������� ��+=OZ�\�R�ht	%c��y �� � �txtP�t  ��R�8�5G>Y� L�^� ������// '/9/K/]/o/B�|�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�/�/�? �?�?�?OO1OCOUO gOyO�O�O�?�?�O�O �O	__-_?_Q_c_u_ �_�_�_�_�O�O�_o o)o;oMo_oqo�o�o �o�o�o�_�_�_% 7I[m��� ����o�o!�3�E� W�i�{�������ÏՏ ������A�S�e� w���������џ��� ���&�O�a�s��� ������ͯ߯��� '�9�4�F�o������� ��ɿۿ����#�5� G�B�T�}Ϗϡϳ��� ��������1�C�U� g�b�tϝ߯������� ��	��-�?�Q�c�u� p߂߂��������� �)�;�M�_�q����� ���������% 7I[m���� ������!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�� �?+?=?O?a?s?�? �?�?�?�?�?�?�/�/ 'O9OKO]OoO�O�O�O �O�O�O�O�O_OO G_Y_k_}_�_�_�_�_ �_�_�_oo_,_Uo goyo�o�o�o�o�o�o �o	-?JcLaBa�Xudy%Sv}�v�y�t� �
�d}xds@cdu  ��Ba8�%�7�>I�� <oNo ��������Ϗ��� �)�;�M�_�2ol��� ����˟ݟ���%� 7�I�[�m��z����� ǯٯ����!�3�E� W�i�{���������տ �����/�A�S�e� wωϛϭϨ������� ��+�=�O�a�s߅� �ߩ߻߶������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ���������1CU gy������ �	?Qcu �������/ /)/$6_/q/�/�/ �/�/�/�/�/??%? 7?2/D/m??�?�?�? �?�?�?�?O!O3OEO WOR?d?�O�O�O�O�O �O�O__/_A_S_e_ `OrOr_�_�_�_�_�_ oo+o=oOoaoso�o �_�_�o�o�o�o '9K]o���o �o�o����#�5� G�Y�k�}�������� ������1�C�U� g�y�����������Ώ ��	��-�?�Q�c�u� ��������ϯ�ܟ� �)�;�M�_�q����� ����˿ݿ����� 7�I�[�m�ϑϣϵ� ���������
��E� W�i�{ߍߟ߱����� ������/�:�<�2��H�T�%C�m�w�ocykd�� me=T�xT�0�T�  ����2�8���'�>9�� ,�>� w��������������� +=O"�\�� ������ '9K]oj|� �����/#/5/ G/Y/k/}/x��/�/ �/�/�/??1?C?U? g?y?�?�?�/�/�?�? �?	OO-O?OQOcOuO �O�O�O�?�?�?�O_ _)_;_M___q_�_�_ �_�_�_�O�Ooo%o 7oIo[omoo�o�o�o �o�o�_�_�_!3E Wi{����� ���o/�A�S�e� w���������я��� ���&�O�a�s��� ������͟ߟ��� '�"�4�]�o������� ��ɯۯ����#�5� G�B�T�}�������ſ ׿�����1�C�U� P�b�bϝϯ������� ��	��-�?�Q�c�u� pςϫ߽�������� �)�;�M�_�q��~� �ߢ���������%� 7�I�[�m�������� ��������!3E Wi{������� ���/ASe w������� //+/=/O/a/s/�/ �/�/�/�/�/�/�� '?9?K?]?o?�?�?�? �?�?�?�?�?�/?5O GOYOkO}O�O�O�O�O��O�O�O__����$PURGE_E?NBL  ,A-A��-A4PW}F<PDO  DT4,BOQ TR_I]TgQ�KUTQRUP_�DELAY ��"A"AKU,B�R_HOOT %�UiR%+B��_�]�SNORMA�L�XKR�_!o�WSE�MI o&oeopQQS�KIP_GRP �1ĞUMQ x 	 ho�o�o �o�o�o�i�U'w GYk1�}�� �����1�C�U� �e���y�����ӏ�� ����-�?�Q��u� c���������͟����)�;��U�$RB�TIF^T�ZY�CV_TMOUT^V�U��Y�DCR�cƾ�i ��a>��0?,AD�v��,ACM�� �����	���,A��=$,A�����o�ȯ ;���;aʤ;�r�@;��;�	�<$D�p/@�j�{� {� ����ſ׿����� 1�C�U�g�����vϯ� �Ͽ�����	�L�-�?� ��c�u߇ߙ߽߫��� ������)�;���_� J��n������ � ��V�7�I�[�m�� ���������������� ��3WB{f� �����*�/ ASew������,kRDIO_T�YPE  �[���REFPOS�1 1Ǟ[
 x	SoY)�}/��/ �-L/^/�/�/�/?�/ A?�/e? ?b?�?6?�? Z?�?~?OO�?�? O aOLO�O O�ODO�OhO �O_�O'_�OK_�Oo_ �__._h_�_�_�_�_ o�_5o�_2okoo�o�*o�oNo�o�o/%2 1�;+J/�o�oL �opvo�/��� ����6��Z�l�-'3 1�
�� V�ԏ��������@� ۏ=�v����5���Y�x�p�0$4 1ʍ� ����۟Y�D�}����� <�ů`�¯��������C�ޯg���0$5 1���&�`�޿ɿ� �&���J��Gπ�π��?���c���z�0$6 1�;+�������`��τ��3!7 1��.�@�z������>��S8 1α��������x��/�SM�ASK 1�� pH ������XNO����4�D�/!MO�TE  �M�_CFG �[�D�."PL_RANGW��+!_���OWER �;%��g�."�SM_DRYPR/G %;*%X� ���TART ����
UME_PR�O����j,$_EX�EC_ENB  y�c�GSPDC ̅ �e��GT3DB��
RM��MT_��T��Y���OBOT_ISOLC����x'NAME ;*�KJLTVL�211350R0�1J_ORD_N_UM ?��
!_H6�8��895  ��+!���������|� ��/ PC_TIME�OUT�� x/ S7232t�1�;%�� LTEA�CH PENDA�N�p�G�I�n�W��Maint�enance C�onso�C�R,"�b/��	UnbenutztY*�/X/�/��/�/�/�/�b"NPqO �K����SCH_LF ����	�1T;MA�VAIL��5���c�SPACE1 {2��
 K?@HHG�v�F�������4L8�?� L;WOL?;O�O�O�O�O �G�?OO%O�OIOkO ]_~_A_�O�_�Y�#� �]�O__%_�_I_k_ ]o~oAo�_�o�o�o�O �_o!o�oEogoYz =�����o�o /�Suw9��� ����������+� ُO�q�c��������� ��ߏ���'�՟K� m�_���3�������˯ ����#�ѯG�i�[� |�?�������ǿ��� ��1�C�U�WϾ�;� �Ϯυ������	�� -���Q�s�e�7߉ߪ��ߓߥ��52�?�?�� �#���G�i�x��\� ����������*�<� N�`�r�t���X����� ������&�8�J��� n����T���� ��"4F�j� ~�R���� 0B�f�z/�/ ^/��/�/�///,/ >/�/b/�/v?�?Z?�? �?�?�???(?:?L? �?p?�?�?VO�O�O�O �O OO$O6OHO�OlO �O�_�O�_�_�_�_�O _ _2_D_�_h_�_|o �oPo�_�o�o�o
oo .o@o�odo�ox�\ ������3��
� .@�d����� y�ˏ�ӏ�5�G� Y�k�}�������u�ǟ 蟿����1�C�U�g� �������q�ï��� ͯ�-�?�Q�c���� ������o����ٿ� )�;�M�_�σ����� ��{�ݿ�����%�7� I�[�	�ϡϓߴ�w� ��������!�3�E�W� i��߯߱�s����� �����/�A�S�e�� �������������� �+�=�O�a����� ��m����' 9K]����@y���/�4� '�9K]/���/ �/�/�/	?�/?#R/ d/v/�/�/�/�??�? �?O�?O<?N?`?r? �?2O�?�?�O�O�O_ _�O8OJO\OnO�O._ �O�O�__�_�_o�_ $oF_X_j_|_*o�_�_ �o�o�o�_�o Bo Tofoxo&�o�o�� �����>Pb t�4������� �ڏ�:�L�^�p��� 0���ȏ���ޟ��� ��6�H�Z�l�~�,��� ğ��ׯ�������"� D�V�h�z�(��������ӿ���	���#+52.D/V�h�z�(Ϟ� �����ϳ��&��;�#+6O�a�sυϗ�E� ���������"�C�*�X�#+7l�~ߐߢߴ� b�����	�*���?�`�G�u�#+8����� ������&G
\�}d�#+G �N5+ �:
�  �,: 5%K]o������ ��o�>d � %/7/I/<j/|/�/�/ ����*�/�+?
/ ;?M?_?q?d/�?�?�? �/�/�/�/?O7O*? [OmOO�O�?�O�O�O��?�?�?O$O6_ `� @> oU� }_�O�_�Ek_9_�_-O o�_�_�_�_loo1o So�ogo�A�a�E�c�o �o!�e�oSe �9k���������L
�_n�@��_MODE  ����S ��]�_Z���_��9�	4�]�D�CWO�RK_AD��{{��F�R  ����b���_INOTVAL��������R_OPTION�̖ ��F�TC�F� ۗ���?���7���V_DATA_GRP 2��H�DU@PJ�y�F� ����G�ʯ���ܯ�  �6�$�F�H�Z���~� ����ؿƿ����2�  �V�D�z�hϞόϮ� ���������
�@�.� d�R�tߚ߈߾߬��� �������*�`�N� ��r��������� ��&��J�8�n�\�~� �������������� 4"DjX��Be� �������q�5 #YG}k��� ����//C/1/ O/U/g/�/�/�/�/�/ �/	?�/??-?c?Q? �?u?�?�?�?�?�?O �?)OOMO;OqO_O�O �O�O�O�O�O�O__ _%_7_m_[_�__�_ �_�_�_�_�_�_3o!o WoEo{oio�o�o�o�o ��o� ��o�oA we������ ���=�+�a�O��� s�������ߏ͏�� '��3�9�K���o��� ��ɟ���۟����� G�5�k�Y���}����� ���ׯ���1��U� C�e�g�y�����ӿ�� ����	��Q�?�u� cϙχϽϫ������� ��o>�b�M�ߕ� ߹ߧ��������� �%�[�I��m��� ���������!��E� 3�i�W�y�{������� ������/e S�w����� ��+O=sa ������/ /9/'/I/K/]/�/�/ �/�/�/�/�/�/�/5?�#?Y?+��$SAF�_DO_PULS�  -��������1t0CA?N_TIME�0}���3���1R ������8�		����
�8����4�4��  ^�OO0OBOTOfO�?��O�O�O�O�O�O�G��1  B2�T�1�1dXQ Q��4}��1�� @ CVT[�0P_z_�\�1�_��WP�U�� {@B�3T i_��_�_oiT D��oAoSoeowo�o �o�o�o�o�o�o�+=OaX^?VNV{py 
�q�p��y�3�1;��o}��4p{}
�t� �Di�0��A�1�z�� ��B�1�q�1�A�1�z�Y�k�}�������  ��������  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v���������@Я�����$��h_ H�Z�l�~�������ƿؿ'�>T�Q���R �7�I�[�m�ϑϣ�Žρ�0�22�@U<�}����$�6�H�Z�
��^�^ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x�������������� ,>Pbt� ��#�����`(:L�2��P+�imih��0�A�B Ѓ�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?OO*O<ONOYG�=X��*`YO�O�O�O �O�O�O__&_8_J_�\_n_�_�_�_�_�ZB��_�V�_i���A��_/m	12345678�r�`!B  �/h�@��jo|o �o�o�o�o�o�o�o q �O#5GYk}� �������� 1�C�T�w������� ��я�����+�=��O�a�s�����V�BH��П�����*� <�N�`�r����������̯ޯ�[�;�j ��&�8�J�\�n����� ����ȿڿ����"�4�F�]�D�_wωϛ� �Ͽ���������+� =�O�a�s߅ߗ�Z��� ��������'�9�K� ]�o��������� ����#�5�G�Y�k� }��������������� 1C�gy� ������	 -?Qcu���Ug`���`�/�/%("C��A��_J   �mH2RqBgb%)
�Pdq#+�?`��R2��/��/�/�/�+pM$ZO���/0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O ?�O�O�O�O�O__ (_:_L_^_p_�_�_�_��_�_�_�_ ooG!��$SCR_GRP� 1����� t ��G! R%	 Ra�Zbkbdd�f%f!�e�kwg�o�o�o(-��a �bD�` D���.qcw�k<�R-2000iB�/210F 56�7890� @tX~� RB21 Op�C#
V06.10 zp�hKa�br#
�u�vZa�fIa�cIa3f!�ahj�a�y	�r�
��.�@�P�?��H��r�r�^g�vN� C��*ZDu�D�d�I��>��\�N���Tva�B3���3�l�B���� Y��� :8�m/�P�  = A�C��-�Dd�hZ`�OG!�o��o�1�.'"��h�p��X�eB��_�B�  ~�ǐ�rvaAL ��  @G 井va@�`ʟ  ?������: 򟨛vaF?@ F�`�%� �I�4�m�X�}����� ǯ��믖i������0��%�7�B�E�گ ��v�����ӿ��п	� ��-��Q�<�u��/�� �c�o����i
����4C#�@㒓� ߘg�Ο@�B�P�1234Ns`׀h���C$A�gRa��㏛cd!%2�rG! ��������2�>�P�� Pv�(|����� Ibp`�t Z`�}�{yi��gϩo�i 7��P�����7uIndepe���nt Axes Qs	����n�f�w ��s�w3i��r��� j|����c��	8���ؙ�/ A��Z��~iϢ� S��/������/�� �F/藦�t/��/� �/�/�/�/?�/?=? (?a?P�:�p?�?�?Z� �?R?O�?'OOKO6O oOZOlO�O�O�O�O�O ����#_f�����k_}_@�_.�Rٺ_\�n�~� o��L$o7o��boto �oUo�o�o�o�o�o��S�����_ ��:��._����� ����������p�$ 6HZߏ���'� ���o�~������ Hohퟀ��#��G� �h�
/��./P/R/d/ ���0�1��U�@� e���v�����ӿ�?�? �����?Q�Ŀu�`� �τϽϨ�������� �;�&�_�
�_m�� F_X_�����_�_�_�_�V�_w�o���� ���o�������+�=�@�a�s���$6xB T����3�� W���,�>�P�b� ���������ΏSe w��:�L�^���� //+/��ܟa/��/ �/6��/Z��/~� ?�� įƯدZ?|/�?�/�? �?�?�?�?�?�?#OO GO6� �VOhOzO@��O 8O�O�O_�O1__A_ g_R_�_v_�_�_�_~ ���_L����Qocouo �2�8�J�8ff��o ��4/Z�Wi8 y���������$SEL_DE�FAULT  ~����P��MIPOWE?RFL  6e.��7�WFDO#�� .��RVENT? 1����,���`L!DUM�_EIP����j�!AF_INEx"�Ə�T!FT��������!�>� ���e�!RP?C_MAINf�H�q�T���x�VIS���G������!TP&�PU����d�I��!
PMON_POROXYJ���e8�����c���f���!�RDM_SRV�⯯�gЯ-�!R�Z�I���h�y�!
�z�M����ih�ſ!RLSYNCƿ��8���!R3OS��8��4 �]��!
CE�MTC�OM^ϲ�kLϩ�!=	r�CONS�ϱ�l����,������� B�g�.ߋ�R߯�v��� ���߾�����?�����RVICE_K�L ?%�� (�%SVCPRG1r���2����3�����4
����52�7���6Z�_���7������8������	9������D����� ��'����O����w ��$����L����t� ��������?�� ��g�����=� ��e���/�� //���W/��/�� -�/��U�/��}�/ ��w������B? �?��?�?�?�?�?�? �?OO?OQO<OuO`O �O�O�O�O�O�O�O_ _;_&___J_�_n_�_ �_�_�_�_o�_%oo Io4o[oojo�o�o�o �o�o�o!E0 iT�x�������M:_DEV ����MC=:����%�~�OL   ���i��!�OUT�`�:�~!�REC 1�d5�L��   �d� 	  �* �- ��(��.����% ����L�����K�����C�
 ��W��:6 ����  _�  ]
�e ��� ��d5�����ҔM�m!
 �瑁� UO7��7�� �:7��Z7����7��7�_� ������M�hz7���W�u]�V� ��^��M�%sM�R�� �� �9�� �1���P��7�P�ՠ7�b7��U� �T7�51C�!�Uy��X���]��eEq�I*0��$� �UfR�E}���*���  k �� �gٯ A)17���ѡ7�r ��� ~�7��M������� ����)�Q+j�]����	 � �� �`�s�)� � 5�q�h�y����J��7��L�7�� ���� [퐃�����M���퟊ �@Q�na���l� I ������� ��Rm���� �`1Ͽ�ѿ����� E������� �lQ�S[J�a�#M�q�������?��K6lL�]���� �+ *7�g �Į�7����K�i�=�������0퐍��K�a����d��E ���RM�-�C�j ���a�A�d���]� 97��\��7�G7������7�������h��BM����VBkP�e� ��  �e+!�S��� �� �P�M��߷�t�J�҄ ��7�x��]�eT�$M�~��
�@Ƞ������ ���������G�Y�k�}����M��� ��>
�a ���h��L]�̠`�t��N �� �1��� ���o� ��� N�7�� �87��7�S�7��џ�T��������
J���2 ��z�V�	��-�?�Q� c�uχϙ�S�e�w�������{�����GZ� ��q��M�EJM��� �����5� � �'L!�� �E�������]� �`�J��&1���T %� ��M�4!�� �a���� �� GE/K O �'7��ɔ��m/ ,m��M��*����� ��U�g� yߋߝ���������� ������������/߼A�S�Mp�6y<w������p�!��?�Ѐ�2�IO ���5y��7�x �ؾqO	)���T �������s7�4�K}�e�B ��A �&��8�O�A���3Km�X  �O��b��� �7� %_+ΐ�� �m����(��L{�5�HW"?�ȁ ���ɹ�_+Z�9_����	@�\P� �>�7��*���]�&Z��(���o=M���_
���) �3 �Y�Mo VT�� �Q7��7��I7������T��̦�0r�`����1UG�o!��o����/SF��J�:�]� �7����k����J7Ԅ�]�1���k���7m�s�]���/^������������	�g�LS	g$A,�0i�G�Y�ß��ş˟���N7a�7�����o��)�q�w�a�޿�OPyC�	�`��������.��#��k�Q��j67r _!w�m�K�]�ǿ�*�ɿϿ�� ���%�K�9�o�]ϓ� �Ϸ��ϫ�������� !�G�5�k�M�_ߡߏ� �߳�������ܒQ�0Ae���	��QT ���q��������� )�OVQ��u�ˏݏ ��e���%�������) ��M;]�q�� ��/�&L�.��17!K}���+ˁ_q�Yd����+/� ;/=/O/�/s/�/�/�/ �/�/?�/'??7?9? K?�?c?�?�?�?�?�? �?�?#OɯۯYO/eO kO5��OyO�O�dL_ H)__M_8_q_�_6� O�O�O�_�_�_o�_ %o7oo[oIoomo�o �o�o�o�o�o�o3 !WE{�o�� �����/��#� e�S���w�����я� ŏ�����+�a�O� ����y�����ߟ͟� ��9��]�K�m��� ������ۯ�ϯ��� 5�#�Y�G�i���q��� �����׿���1��L �_,�v�dϚψϾϬ� ��������$�*�<� r�`ߖ�xߊ��ߺ��� ���� �J�,�n�\� ~������������ "��F�4�j�X�z��� ������������ BT6xf��� ����P >tb����� ��///L/./@/ �/p/�/�/�/�/�/D� n_'??K?6?o?Z?�? �_X��/ ?�?�?�? O ODOVO8OzOhO�O�O �O�O�O�O�O�O.__ R_@_v_d_�_�_�_�_ �_�_�_�_*ooNo0o Bo�oro�o�o�o�o�o �o&68J� n������� "��2�X�:�d�j�|� ����֏ď����0� �T�B�`�f�x����� ����ҟ���,��P� Fϸ?^�`�������� ί����:�(�^�L� n�p����������ܿ � �6�$�Z�l�Nϐ� ~ϜϢϴ�������� �D�2�h�Vߌ�zߘ� �ߤ���������
�@� .�d�v�X����� ���������$�*�<� r�`������������� �� &8nP ~�������f��$SERV_�RV 1�	8��0(	\�n���!3TOP1�0 1�=
 �6 q�. 2V#Tq� sE� q�6r _�*$�*" *q�� E�YPE s q��H�q�1HELL_CFG �t&�0��? �?�/q�%RSR�/�/�/? ?:?%?^?I?�?m?? �?�?�?�? O�?$O5M�DD<I�  �E%5OvO�OCE?Mbq��O�B�@�D�\D!d�Oq��)�}&HK 1�+ P"�O?_:_L_^_�_�_ �_�_�_�_�_�_oo�$o6o_oZolo~oz)OMM �/�o|"�FTOV_ENB�i$Et*OW_RE�G_UI�o{"IM/WAIT�b�I{�OU! tDyT�IMu��WV�AL,s_UNIaT�c�vt%QLCpWTRYwt%1�MB_HDDN �2�k P  �����>�5�G��t�k�}�����̌�qO�N_ALIAS k?e�iLhep� ��(�:�L�D��w� ������X�џ���� �ğ=�O�a�s���0� ����ͯ߯񯜯�'� 9�K���\��������� b�ۿ����#�οG� Y�k�}Ϗ�:ϳ����� ���Ϧ��1�C�U� � yߋߝ߯���l����� 	��-���Q�c�u�� ��D���������� )�;�M�_�
������� ����v���%7 ��[m��N� ����!3EW i������ �////A/�e/w/ �/�/F/�/�/�/�/? �/+?=?O?a?s??�? �?�?�?�?�?OO'O 9OKO�?oO�O�O�OPO �O�O�O�O_�O5_G_ Y_k_}_(_�_�_�_�_ �_�_oo1oCo�_To yo�o�o�oZo�o�o�o 	�o?Qcu� 2������� )�;�M��q������� ��d�ݏ���%�Ѓ��$SMON_D�EFPRO ����N�� *SYSoTEM*Ё�>��RECALL ?�}N� ( �}�׏����ԟ���  ���/�A�S�e�w�
� ������ѯ������ +�=�O�a�s������ ��Ϳ߿񿄿�'�9� K�]�o�ϓϥϷ��� ���π��#�5�G�Y� k��Ϗߡ߳������� |����1�C�U�g�y� ������������ �-�?�Q�c�u���� ������������) ;M_q��� ����%7I [m ����� �~/!/3/E/W/i/ �z/�/�/�/�/�/�/ �/?/?A?S?e?w?
? �?�?�?�?�?�?�?O +O=OOOaOsOO�O�O �O�O�O�O�O_'_9_ K_]_o__�_�_�_�_ �_�_�_o#o5oGoYo ko�_�o�o�o�o�o�o |o�o1CUgy ������� �-�?�Q�c�u���� ����Ϗ�󏆏�)� ;�M�_�q�������� ˟ݟ��%�7�I� [�m� �������ǯٯ �~��!�3�E�W�i� ��z�����ÿտ��� ���/�A�S�e�w�
� �ϭϿ������ψ���+�=�O�a�s���$�SNPX_ASG 1�������� P �0 '%R[1]@1.1zߖ �?��%����<��Q����_*_8�G�ֶo�6�w�� �.�f��֦�8���� ׯ�#������ ���7��$��E&�g���K8V���֟8�����֡0������!��0��'� t�W��� ��� �v��/q����v���
�2G
�1�6w����� ׆��� �l1G�/����6/� �Q�&/g/�Qc<V/�/����D�/h	�/�/ ��/&? ׄ��?W?I�qF?�?�&�v?�?�2�Y�?�?���ϴ�?O�׋8OGO���6OwO���?�OY�|x8�O�O�	�O_��n�M�O7_��c	�&_g_��߅/�_ �J�\�_�_�c�5O�_ ��u?�&o��5OoWo�Oq�Eo�o �]o�vo��o�獦o�o�z1b�� �ޒ%/F� יC�Ov����f�:� ��7q�/� ������7��'AJ&�g�ֵq��� ע�%��ǏւA/�������4��'��~1j�W��@���� ��I�v�����>1w���ZwN�֟���R�u�F� ���1�6�w��'�f����֑����ׯ��16�O� א��6�"�I|&�g� �'��p�ߋ�̿Ѹ����� ��'Ϫ��]ώ��#tFχ�և���R��PARAM� ���� �	�P<�P!�I��D���OFT_K�B_CFG  �]��ԉ�OPIN_�SIM  �����=�O�a�Q ��RV�QSTP_DSB�&����h��SR� �)� � �& FOLGE�124 .����0�022A��Ī�TH�I_CHANGE7  �E��GRPNUM� ��OP_ON_�ERR��I�PT�N )���C�RING�_PR1�U���V;DT+� 1�ɑ@�@���F�������� � �1�C�U�g�y��� ������������	 -?Qcu��� ����); M_r����� ��//%/8/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_P_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�h�y��� ������ӏ���	�� .�?�Q�c�u�����e��VPRG_COUNT��|��ƒ'ENB����M�4�~��UPD 1���T  
����B� T�f���������ׯү �����,�>�g�b� t���������ο��� ��?�:�L�^χς� �Ϧ����������� $�6�_�Z�l�~ߧߢ� �����������7�2� D�V��z������� �����
��.�W�R� d�v������������� ��/*<Nwr ������ &OJ\n����������_CTRL_NUMГ�!�!"GUN�%" 2�0�� C 1$4!!4!/s$A
1$Ւ(#�'�/�/�/�/ÐYSDE�BUGА1�� d��� SP_PAS�SЕB?;LOoG �0��� J1�^���k$[=�%UD�1:\04.12_MPC6? c(�?g=�x82�?�2SAV� �9=�!n%&�x8SV�;TEM�_TIME 1��R+ ( @���"1��&���#hF�sO�O�L�٧O�O�O �T1SeVG S+�ѕ'���PASK_OPTIONА0��ߑ'Q_DI0�ߔ�TBCCFG ��R+�=�.�_`�_���!�_�_�_o �_5o oYoDo}oho�o �o�o�o�o�o�o
 C.@yd���@���	��%� 6��i�{��X����� Տ�����0��=P� !�G�5�k�Y���}��� ��ßşן���1�� U�C�y�g�������ӯ ������	�+�-�?� u�[�F�������˿ݿ [����7�%�[�m� �Mϣϑ��ϵ����� �����E�3�i�Wߍ� {߱ߟ���������� /��S�A�c�e�w�� ��������+�=� ��a�O�q��������� ������'K9 []o����� ��!G5kY �}�����/ �1/��I/[/y/�/�/ /�/�/�/�/�/?-? ???c?Q?�?u?�?�? �?�?�?O�?)OOMO ;OqO_O�O�O�O�O�O �O�O__#_%_7_m_ [_�_G/�_�_�_�_�_ {_!oo1oWoEo{o�o �omo�o�o�o�o�o /eS�w� ������+�� O�=�s�a�������͏ ���_	��9�K�]� ۏ��o�������۟� ��͟#��G�5�k�Y� {�}���ů���ׯ� ��1��A�g�U���y� ����ӿ������-� �Q��i�{ϙϫϽ� ;���������;�M� _�-߃�qߧߕ��߹� ������%��I�7�m� [����������� ���3�!�C�E�W��� {���g������� ��A/Qwe���� �$TBCSG_GRP 2����  ��  
 ?ú�����  <N8r\ ������� �/,//P/:/t/�/ l/�/�/�/�/�/?�/ (?:?$?^?D?n?�?~? �?�?�?�?�?O�?6O�HMA��*SYS�TEM*� V8.�2306 qC4/�2x@014 A� t  _F_GF��� PARAM_�T   ��$MC_MAX_�TRQ��$�D_�MGN�CC� AV��ISTAL�IBR�K�INOLD�FS�HORTMO_L#IM	Z�M�EJPTWPL1CU2CU3CUU4CU5CU6CU7CU8�A `�A��A�� �_ACCEJR�WTQ�SPATH�W�Q�S�Q?_RATIO�B�S��@ 2  	$�CNT_SCAL�E	ZSCL�CIN^�Q_UCA��b�CAT_UM%hY�C_ID 	*cB`_EKPGjTPGj�]PG`PAYLOA�WJ2L_UPRo_ANG�fLW�k��a�i�a�ER_F2�LSHRT�gLO��da�g)c�g)cACRL_Shpgzd�BHVA`  �$H�B:rFLE-X7s<�@Jb�@� :$aL�ENKQguTQ$DEjx�t|s�R�X�p��zSLOW_AX�Iq$F1aI��s2�x1�q�u�wMOVE_TIMd_INERTI%`�:p	$D	�TOR�QUE�Q!��p�I>HPACEMN�`�(�P�s�E^�V�p�Ap/�x�@�x�TCV����@��A�������@T".��@��J�Aꉄ���M	�(a�(`J�_MODa�p�S R�@�gq2�@	P�^�Eo�0`J�遉Xp�A�RU�?�J�K.�����KKSVKvTSVK]SJJ0딶KSJJTSJJ]SAmAKSAATSAA
�ffSAAoS�AN1ǌ�<����@�@PE_N�UQ� VqCF�G�A � $�GROUP�@SK�&cB_CONFL�IC�dB_REQ�UIRE.q�qBU� sUPDAT�v� �ELk�� Τ�^�$TJ�P�;JE�@CTRa�q�TN	�F˦��HA_ND_VB8rVq�OP�U $]�F�2�F
�TSCOMP�_SW&a�@�@�F?� $$M�`�IR�C|��A��x��R&��A_}b�FDļ�MUA�LA�LA�KA [TҰ�KD�LD�KD [�P�PGR�Gp�ST��Gp��Ip�NXDY�`R�@�E��ڵ�` ` �g�q�g�a�g0�<Q@��p��UPKUTU]UfU0oUxU�U�R Vr�T� r�Wt�R �%�n�TPy�ASYM$�U:p� �V�Pm�ao_SHo�g4d ]��C�>oPoboto�cJ�l>P�j^�T�i
�_VI&���Ѫ�V_UNI�c��TS�aJ��������l�� �e����m�y>P�1a���GtOsq����TCPPIR�A  ��ENA�BL�p����$T�CDELAYݱ�
��SPEE4P ? X ��I�!N� ސ��� GP��`��Q���q�@MPڢ�PROG_���Y�PEڡ��_z�	 1|�m���SE s���m���' ǦWARN�I��EN&���OT1F�qj��_T���SMAARSCW�t��wSPDz�
 �������EARTBE����ET��z���P�PARGAT��FLQG�u�|sS�@E�@R&�6�%�aos6REAJVXTR܉� OUT�A !p렜��� E��̢�ID`�(d^�U c�A�`��޵�G��Q# �PH����<��{I�$DOp����z� �
�I��A��J �p���W#�۠�� ���� � T�MEJS���R���T EP��"@Pl���#��(�!�)T"�m�� $DUMMY}1]Q$PS_�p�RF�pg@$�&��FLA|��2�GLB_Tu�k*5����(���8!������QSTT���SBR�PM21�_V�T$SV_�ER�`O�p3�3C�LD0p2A^����G�L��EW�A 4l��$��$Zݲ!W�3���`P�As %b� �3U�5 �]�N�0�$G�I�}$�1 ���1�0�A L���F�}$F�ERFN� M�NcF]I�J�TANCb��J� RǱ �1$�JOINT����$I0�1M� �Q��FECE�q��S�b��*B|���Q� �p�US�?��LOC�K_FO�`[�� B�GLV��GLXT�  _XM`�AEM�P�@�� -PB2�@G$US�!�0p2*��4QQRW��@QQ��SCEj�CrP $�K��M#TPD�RA�0�T�AVECXlp�V�@IUQQVQ{HE�@TOOL�s��SV�tRE�PIS�3|s�T64�)`ACiH� ���QON���$29�"�PI� � @$RAIL__BOXE���oROBO"T?�r1�HOWc>d� aROLM�"ge_�
dxbp��/`�p6�O_F��?!  
�2�QR^q�N��R�PO]ra�B�p�A�`ģE~X2MU�֡��,�@	 IP#VNK��R�/b�Q
�QQ�`�PCORDED�@���`�A���OY   D )0OB�٣�@�dwSq�#E Sr�ۡS;YSSqADR =Q�TCH��  �, �A�A_D��th��A'AVWV}A�� � �P��2kPREV_R�T��$EDIT��VSHWR��p��$�K��IND� R`;�$��D&�h[�U�6��KE��� �l�JMPppL�jX�TRACE�)[p�I,PSڢC �NE�Pۡ��OTICK�S��Mo��t��HNR1 1@]p��L	_GK&fΩ�STY�aLO�D1�b����~� �t 

 G�u%$��qD=� SFp!�$��8��!�F �P���LSQUaLyO���TERC� �ݱ��Sz�  @h0�� p��㡼Q,�1O� �#dIZ4A��! C�"!�o�UTPU��1�_DYObB�pXS�@Kj�AXIP��cVQU1R���0i#$TH`��~vK���_�P�rET���P Rlp��O�Fd��P�A�����$� cc>   �qS=R3� lѐu� �a����������� �ù�ӹR���R�� R��d�~�B�d�������C翐�C��� �2�D��SSC,0 o! h�0DS�4� X}�AT��<��� ~���"ADDR�ES�SB�SHIyF�HP_2CH�p�zqIK0���TX_SCREEUr"	 =k�TINA�3@���D�1����T0# T���0'�g00��^��r^��RRO�R_vA��(�h$�UE5$$ ��Щq09S�1�qRSM��T�UNEX��j���S_�3��G�ѽ����G�C�B��� �1#�`UE�%�="�2��MT!�L�v�m�w0O�D\��UI_� HP� O& 8e�w@_T���f� R���Bcg��" �R�O��T0'����7$BUT�T��R RraLUM���u���ERV��R�Pa@��S1({ ^ƠGEUR&SF����A)� LP���E��C�)#�S�1�c�1�T�P0�5.�6.�7.�8����a@����%�Q�AS�'�R�USR�4) I<Z0� UB�AI΀�@FOC�Q@PR�IΡm`�� TR�IP�m�UN$ 5$*	@t�$ k�cj�HR���� �+a��� �G `\��1���\OS��qR��V�H�QS1,��?�3�>���`HRU�S1-������NHOFF!PT0.[p��O' 1,�09-�0GUN?_WIDTH�b�B_SUB�"p0�'SRT� �/��vA̗` �OR`�RA�U��T����VsCC�М�0 �aC36MFB124��VC/0.D1h# %bTq���4.Ȕ�c)�C�`	%DRkIV���_Vu��,$(��@D��MY_UBY��$V�vA��  B�tC�#�QtBi0pp�+��"L7�BM�1�$��DEY!�EXpG�n��Q_MU��AX�10orbҲ�Gð�PACIN΁}�RGC�52�2�32���!RE{����Q�b��2�02�TARG�@P1Rc0�`r�R� �03 d��N_�FLA΀r	�"�N�RE�#SW0_AA1�`�@�!�O���A���3�E��U�B�a�`���HKG�4���:�����05�!CEA��+GW�OR!P�5
�4MR�CV�5 ���O*S�M!PC2S	hB`3hBREFF�FqF \A�0�࿣�0��mJ�A�~J�A�K�EqFO_R!C,KXEKV�S���'�]#�q�5�6 �$���1؄��b%�p�ROU�[2�# �1z52�2�P$0���� �΀3��2����Kq�SUL��14;r��6�5� �P @�3�cN�f��f��c�PL�#5e�#5e���Ag���$��7G0 &��ǡ4� ��C�`+�LO�A�d�a�� �iu��`ܓC�pM-I��FR�hTj��fNR[$HOh��r�`�COMM'#��OB��v{X���؇VPx]2�Hq_SZ3c2Qu6/cQu12��Nx�0Lx�`LxWA�eM]P�zFAI�`GT��`AD�y�!IM�RE~T�r_�GP��� ��&ASYN�BUF�&VRTD����qσOL��D�_�:�W�P�E�TU�#�`Q�0�EwCCUP8VEM:0x�e���gVIRC�q�2�`le�8u��0C�KLAS^	�V�LEX��9/d�����	�LDLDE�FI<� �r�.������Tp�Q���:����Tp1�'�����V�� ;`��L���{,f�"UR�3�0_R�p 󔟑�!���U3�/�/��$�`7���0Ғ �T9I�Q��SCO�� �Cz�4;#6;�; �;!�;/�//%*�ᢕ���D�SЧ@� �SM<�)���J*��%�ģq�=)G�eLI�N���W�@XSGAq�>  ��N�BPuK�cH��HOL��{&�ZABC}�?v2`�XS�@
�Z/MPCF}@<���2?��l!LNI��@�
t��� ~A ����q+@��CMCM�0CKsCART_�ٱ�DP_�� $J����������S��S��BUXW� ��UXE�!A�<��9��d�J�\�J�~l� (�ZPץ!B���RR�^���uY!�D" Ca�:���IGH&3G�#?(!�!��A@��>�D � T��A�~�$B�PK�'3PK�_a�	c�RV�`F8��Ba�OVCY��@��TU�O0��j�
R�I��1uD��TRA�CEx�V
1��SP�HER��E ,�!��������$T�b� 2������ �d ��?� �	 HD)uˀ� (�[5�0��A��(�$�B����O�Z�$�333.x���<�|Z�\�&�8�������C���� CA?��Cp������θ�|EP��Gz�2�6���sz����	z���@����� ������&C n��p��	�V3.00�	�rb21�	*�� ����
fffjtU�Tp	 ��   ?���Cz�_f�x�� �� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?O��	 O2OO ^OlI0pO�ODlO�O �Kz�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>PbO>O �JO���O��O� (��O0�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯t� ��.��B��v�舿���J�� v��  f+���2f�##���	2?� *�c�Nχ�rϫϖϻ� �������)��M�8� q�\�nߧߒ��߶��� �����#�I�4�m�X� ��|���������� ����8�#�\�G��� k��������������� "XC|�� �I�s�����! E3UWi�� ������/A/ //e/S/�/w/�/�/�/ �/�/?�/+??O?a? k��p?�?�?>?�?�? �?�?�?OOBO0OfO xO�O�OZO�O�O�O�O �O_,_>_�O
_t_b_ �_�_�_�_�_�_�_o o:o(o^oLo�opo�o �o�o�o�o �o$ H6X~l��� ����?�&��?� h�V���z�������� ԏ
��.����d�R� ��v�����П⟜�� ����*�`�N���r� ����̯��ܯ��&� �J�8�n�\�~����� ȿ���ڿ���4�"� D�j�Xώ��:����� tϢ�����0��T�B� x�fߜ߮����ߐ��� �����P�b�t�� @����������� ��L�:�p�^����� ���������� 6 $ZHjl~�� ���� 2��J \n����� ��/
/@/R/d/v/ 4/�/�/�/�/�/�/? ?�/<?*?L?r?`?�? �?�?�?�?�?�?�?O 8O&O\OJO�OnO�O�O �O�O�O�O�O"__F_ 4_V_X_j_�_�_�_�_ p�_ o�_�_Bo0ofo To�oxo�o�o�o�o�o �o,<bP� ���v���� (��8�^�L���p��� ��ʏ��ڏ܏�$�� H�6�l�Z���~���Ɵ ���؟���2� �B� h�o������N�ԯ¯ ����.��R�@�v� ������j�п����� �*�<�N��^�`�r� �ϖ��Ϻ������� $�J�8�n�\ߒ߀߶� �����������4�"� X�F�|�j������ �������$�6���V� x�f������������� ��,>��NPbp����  � �� �����$TBJOP_G�RP 2���� ?���C�	�E�� �����X���y�^ ��,X� �@� ?���D�)̴C2
�C랔���R;#��8����>��$�k<�p�S�>�B��?T�?B��B��rB6�� �'/2'���j/|%�<?D!?���?L�#C  B�Z'�/:/L/^/�/�4[5�2A���;�ŗ-C0�hB�h�/Q?C�d6���Cw�p��.|E�6��?�'�;���C�A�?-�N?�a��1C��xC+9R?�?d?v?�6x4O�6;�?y)�2 ?Gu�PA�CeykC#CK �?qO�?O B�E�O7K�l��2333?_fff?Y-Z�@rO�O�;�%_�'4_ _,_Z_�_f_ _�_�_ �_�_�_o�_�_:oTo�>oLozo�o~D����� ��%	V3.�001rb21�*�`��w� F�� F��. G
� G�(� GG� G�gs G�� G��v G�^ G����G�@�G��; G쑀G��C�H	(�H�� H��H�&��H1�H�;y� r?� F�M4 Fj0 F��` F�v F��V F� G�> G7� G�Zj G�l G����G���G��� G�� G����HS@H���H0) H�B�@=� <��U��l:� R� Z@jQ����
�?�  ��oK�y�� `�\�n���� G����ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �ߪ y���߬߮ !p ���(�:���^�p�� ����	������ j�)�����u�?��� ���������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O���߳O��S��O_ _�O�OK_]_o_�_�_ �_��_����_1�Y� #og�y�ko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i��O�O���O7_ տ�����Ϳ/�A�S� e�wω��_���_�_������$TCPPACTSW  e����IR� e����CH%�SP�EED 2� �C�e�  U�����_CFG %	2�?Ѵ���!�z���_SPD�ӱ
�>Ѵ�<?�:�o���������NUMд���
~��OUT 2��
  ����t��n� ������������� /�"�S�F�X�j�|���ZERO��  ����ESTPARaS�?����HR��ABLE 1��I�Ҋ��ٔ���E�����Ѯ���	��
����⊔�����4���RDI��<�&8J\�O��� �0��S��� �
�//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?�� ���z�w���Y k}�����n2/� 2�P`�0 03�4����2�A�@��`�IMEBF_TT���5�զ��CVER2�!ѯF��ޜ@R 1�8�ﴰ� W cm��7a�6��լ�O����PP�\�$_hY�D�P��0[�\_�[Q�R[Ĕ_�_�_Ř�_�_�_�oGh��Lx���HB[Ǭ�DooX�<o~Niݬx�`o��to�i�t	ݛ �o��oE	B�oVˬo�
;SI�T��inX͌Lf���~�n�rV����S_E�"V�4��oX�}�o�d���]Ҥ�����2V�܏F�T_��������93�3�E����1h�z���� �q�������������uc?��"���_[/�Y�k�'���������*B��ί����������g�9�K�ǉ�`�r�L�w@������D.�!�@��� �MI_CHA�N�G 
�DBGL�VL�G���ET�HERAD ?j��i����0r��:eu�4:34:�2e:91 r�2(��5���4P�RP��@!��!�����~�SNMASK^����o�255.�$�0��#�5�G߁�O�OLOFS_DI����L�ORQCT�RL �ɦ3�:��5�T������� �0�B�T�f�x��� ���������������;�*�_���PE_D�ETAI<ȉָAP�GL_CONFI�G WIgA�?�/cell/$�CID$/grp1c�?�c����������2(]o ���4��3��@�)���40 ew���<��� ��/ /2/�V/h/ z/�/�/�/?/�/�/�/ 
??.?�/�/d?v?�? �?�?�?���}S?�?�OO*O<ONO  O�uOTN�R?�O�O�O �O�O_L?)_;_M___ q_�__�_�_�_�_�_ oo�_7oIo[omoo �o o�o�o�o�o�o �o3EWi{�� .������� A�S�e�w�����*��� я�����+���O� a�s�������8�͟ߟ ���'���K�]�o�������������User Vie�w ��}}1234567890� ����0�B�J�Ӱ��j���ΩK	�?����Ͽ��� e�w�բ �	��_�qσϕϧϹ� �*ψ�SN��%�7�@I�[�m����ψ�5�� ����������u�7�}�6��p�������)���}�7_�$�6��H�Z�l�~����}�8 ������� 2���SY l?Camera٪����������BE �.@�Zl~0�����  r�� �//(/:/L/^/ �/�/�/��/�/�/ ??$?K�rBɻ/p? �?�?�?�?�?q/�? O O]?6OHOZOlO~O�O 7?I7��'O�O�O __ $_6_�?Z_l_~_�O�_ �_�_�_�_�_�OI7� �_Jo\ono�o�o�oK_ �o�o�o7o"4F Xjos^��o�� �����o2�D�V� �z�������ԏ{ I7�k� �2�D�V�h� z�!��������� 
��.�@��I7��ן ������¯ԯ母�
� �.�y�R�d�v�������S�e�98����� #�5�G��X�}Ϗ�6� �����������߮�	t0��Z�l�~ߐ� �ߴ�[������ߣ� � 2�D�V�h�z�!�3�y  {�������	��-� ��Q�c�u�������� ��������t���? Qcu��@��� �,);M_ @�S;����� �/�)/;/M/�q/ �/�/�/�/�/r��K b/?)?;?M?_?q?/ �?�?�??�?�?OO %O7O�/�+k�?�O�O �O�O�O�O�?__%_ pOI_[_m__�_�_JO ��{:_�_oo%o7o Io�Omoo�o�_�o�o��o�o�o�]  �Y>Pbt���������  � y?���B � *��]>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V��h�z�(x  
�`(�  �2p( 	 �������ο� �(��8�:�Lς�p�Цϔ��ϐ�z �^o�!�3ߦoW�i� {ߍߟ߱߸S������ ��F�#�5�G�Y�k�}� �ߡ���������� �1�C���g�y����� ����������	P�b� ?Qc������ ��()pM _q������ �6/%/7/I/[/m/ ���/�/�//�/�/ ?!?3?E?�/i?{?�? �/�?�?�?�?�?OR? /OAOSO�?wO�O�O�O �O�OO*O__+_rO O_a_s_�_�_�_�O�_ �_�_8_o'o9oKo]o oo�_�o�o�o�_�o�o �o#5|o�ok} ��o������ T1�C�U��y����� ����ӏ���	��b� ?�Q�c�u���������@ ��ȟڟ쟻������)fr�h:\tpgl\�robots\r�2000ix&�b�_210f.xml��P�b�t�������`��ί���� �dummy"�;�?� Q�c�u���������Ͽ ��
��.�;�M�_� qσϕϧϹ������� ��*�7�I�[�m�߀�ߣߵ��������� ���)�;�M�_�q�� ������������� %�7�I�[�m������ ����������!3 EWi{���� ����/AS ew������:�;� �88�?�� "/�/@/B/T/v/�/ �/�/�/�/�/?�/? B?,?N?x?b?�?�?�;��$TPGL_O�UTPUT |��  ?O���3;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_�_�_�_�3 �@2�345678901�_�_�_�_o o(c ��_Ooaoso�o�o�o Ao�o�o�o'�o�5]o���=�}�����%�� �[�m��������M� Ï����!�3�ˏA� i�{�������I�[�� ����/�A�ٟO�w� ��������W�ͯ��� �+�=�կ�s����� ����Ϳe�ۿ��'� 9�K��YρϓϥϷ� ��a�s����#�5�G� Y���gߏߡ߳�����?}}!��+�=�O�a�r�@/���*? ( 	 �_�� �����%��I�7�Y� [�m������������� ��E3iW� {������/�V� "7ew S������RP 
//�@/R/0/v/�/ ��/�/`/�/�/�/�/ *?<?�/`?r??�?�? �?�?�?H?�?O�?O JO\O:O�O�O�?�O�O jO�O�O�O"_4_�O _ j_|__�_�_�_�_�_ R_oo�_BoTo2odo �o�_o�o�oto�o �o,>�obt� ����J\�(� �L�^�<�������� ʏl�ڏ �ޏ��6�H� ��l�~� �������؟ �T��� ��V�h� F������¯ԯv��� 
��.�@���,�v����*��������������$TPOFF_L�IM K|�ӱ��|��N_�SV�  x��%� �P_MON7 CG�*��|�2x��STRT?CHK CE���M�VTCOM�PAT:���I�VW�VAR Z�,��h��� ��|��m��_DEFPROG %���%FOLGE1�2��Y�t�_DIS�PLAY���/�I�NST_MSK � �� k�IN�USER��-�LC�K�܊�QUICK�MEN��q�SCR�E�C��t_scq���!�&��%�7�ST��E�RA�CE_CFG UZ����	��
?���HNL �2��#����  ��������"�4�F��X�j���ITEM �2�� �%$�12345678�90����  =<��������  !�����Jӫ� k�����); _�/U�� ��	�7�	/ /?/���A/� �/�/�/3/�/W/i/{/ �/M?�/q?�?�/�?? ?�?A?Oe?%O7O�? MO�?O�O�?�OO�O �O�OaO	_�O�O�O#_ �Oy_�_�__�_9_K_ ]_�_�_�_Soeo�_qo �_�_�o#o�oGo }o/�o�o|�o��o ��SCUg�� ��[��������� -�?���c��5�G��� S�Ϗ��w�ş)�� ��_������^���y� ݟ�����ů7���� m�-���=�c�u�ٯ�� ���!���E���)� ��Mϱ�ÿտY�q�� ����A���e�w�@ߛ� [߿�ߑ��ϧ��+ߔ�߀�S����F�ψ  u�F� 8��P�F�
 ]���j��(�UD1:�\�����R_G�RP 1 ��?� 	 @P��� ���1��U�C�y�g�������s������<����?�  ) I7m[�� �����3!0WEg�	�ա �q��m�/�'// 7/]/���/���/���/ �k�/#??G?5? k?Y?�?}?�?�?�?�? �?O�?1OOAO�� �O��Oe/�O�O�O	_ �O-_k/Q_�/x_�/u_ �_QO�_MO�_�_oo 'oMo;oqo_o�o�o�o �o�o�o�o7uO Se#_�_��� ���M_3��_Z��_ ~��_����ՏÏ�� ���A�/�Q�S�e� ���������џ�E�o5�G��SCB ;2!� ���� ������ϯ�������X_SCREE�N 1"��
 �}ipnl/X�gen.htm$��w���������P��Panel se�tupü}	index.STMÿ���1�C�U�̷
R�obot Info e�9�ϱ��������� �τ�1� C�U�g�yߋ�߯�&� ������	��-�߶� c�u�����4�b� X���)�;�M�_��� ������������� x���7I[m� 6,���!�3�W3�UALR�M_MSG ?D��Q� RD� �����/
// :/@/q/d/�/�/�/m�SEV  {��&kECFG ;$e�  D7�}A1   B�NW�Q�0�4��  A "�X��z2?!�F0�~J?#�Xb?�"NX��z?"�X��?#ز�03�?�1�\�?!UƦ0��?!�1��?�#�0�S�!GRPw 2%e� 0*0�r2�I��I�?2������n��g"6+�,��&0v��O�n��O�O�O�OjI_?DEFPROw+F�� (%FO�LGE124 .�(_-Q0045  �%MAKRO050�OD%�/_j_ �_�_�_�_�_�_o!o�oEo�GINUSE�R  ]�ONoI�_MENHIST� 1&e�  �( P��-/�SOFTPART�/GENLINK�?current�=editpag;e,T5,1�o&D�.�o�o Q011,2N_���9{'HZumenu�b71�o��&�08����a37����������Cq(P�b�8�q24,3u�$�p6�ŏ׏�{190u� v�������E�GYU,1���,�>�I�ߟ�{93�a�o������Ю�6a�a6o��� � 2�D�V�Փ므����� ��ȿڿi����"�4� F�X��|ώϠϲ��� ��e�w���0�B�T� f��ϊߜ߮������� s���,�>�P�b��� ����������ݯ �(�:�L�^�p����� ���������� ��$ 6HZl~�� �����2D Vhz���� ��
/�./@/R/d/ v/�/�/)/�/�/�/�/ ??�<?N?`?r?�? �?�?�/�?�?�?OO &O�?JO\OnO�O�O�O 3O�O�O�O�O_"_4_ �OX_j_|_�_�_�_A_ �_�_�_oo0o�_To foxo�o�o�o�oOo�o �o,>)?�ot ������o�� �(�:�L��p����� ����ʏY�k� ��$� 6�H�Z��~������� Ɵ؟g���� �2�D� V����������¯ԯ �u�
��.�@�R�d��Oz�$UI_PA�NEDATA 1�(������  	�}�/frh/cg�tp/doubd�ev1.stm �8981&action=100p��޿���)prsim�<�  }?��c�uχϙϫϽ� ) ���������+�=�$� a�H߅ߗ�~߻ߢ���������Lv���    <� s�M�/k�arel/pee�ritp ��=1533¿r�����dual����O�  ��$�6�H�Z��~� e������������� ��2V=z�s��#�5� 7ӣ�D���ਸ਼t��3����0B� hirdS}�� ������// C/U/</y/`/�/�/�/ �/�/�/�/?-??Q?�� 4� �$X��?�?�?�?�? �?4?�?O�;OMO_O qO�O�O�?�O�O�O�O �O_�O7_I_0_m_T_ �_�_�_�_�_�_�_p2f��1O6oHoZolo ~o�o�_�o'O�o�o�o  2�oVhO� s�����
�� .�@�'�d�K�����o oЏ����*�}� N��or���������̟ ޟE���&��J�\� C���g�������گ�� �����4�����j�|� ������Ŀ����m� �0�B�T�f�x�߿�� �����Ϲ������,� �P�7�t߆�mߪߑ� ��A�S���(�:�L� ^�p��ߔ�ϸ����� �� ��y�6�H�/�l� S���������������  D+hz��������� )�7��&cu ����$��/ ��;/"/_/F/�/�/ |/�/�/�/�/�/?��������$UI_P�OSTYPE  ���� �	 ?v?E2QU�ICKMEN  �T;c?y?G0RE�STORE 1)���  '�?���?�3�?��mODOVOhOzO �O/O�O�O�O�O�O�O _._@_R_d_Oq_�_ �__�_�_�_oo�_ <oNo`oro�o�o9o�o �o�o�o�_!3 �on����Y� ���"��F�X�j� |���9C�����1�� ��0�B�T���x��� ������c������ ,�׏9�K�]�ϟ���� ��ί௃���(�:� L�^����������ʿބ7SCRE�0?��=u1sc��0u2�3�4��5�6�7�8<�E2USER�쿦��ks�f�3f�4�f�5f�6f�7f�8�f�E0NDO_CFG *T;� �E0PDATE P���KS_2�4�1G�_INFO� 1+�����10�%  OLGE0311п�  �5� G�*�k�}�`ߡ߄��� �ߺ������1��U��g�9��OFFSE/T .�=q�l� �0s����������� !�N�E�W���[����� ��������/y��?{
j���t��SEUFRAME�  d�����R�TOL_ABRT8����ENB��?GRP 1/�9�1Cz  A�: 8l�8J\n��!���
�0U��~�MSK  ����	N�%��%xKH/�2VCCM�³0��]"MR 2=6T9 d�����	��O�~XC56 *�/�&X����0�5��A�@�p��L. 	j8?d�7?I?�v?�!q?�?5�A��l��?�?l�� B����1l��5�?O b??OOcONO�OrO�O �O�O�O8O�O___ M_ Oq_�_d��!�!�/ �_�/�/�/??'?o �O\oSo1_�o�o�?�? �o�?__�o"io{o= jU�y���- ���	�B�U_f�x� ����!�_���_�_�_ oo'o��\�S�1� �����o�oڟ�o_��� "�i�{�=�j�U���y� ����֯-���ɯ�	� B�U�f�x����=��� ��͏ߏ���'�� �\�S�1��ϤϷ�ɟ ���_���"�i�{�=� j�Uߎ�y߲ߝ���-� �����	�B�U�f�x��O/ISIONTM�OU� $r%����d#7�K ��LT/ F�R:\��\DAT�A\�� �� wMC��LOG��   UD1���EX��' ?B@ ��O� ��7/m� �q���� ��  =	 �1- n6  G-��T�L�&,��<���=�����T����TRAIAN6������"8�+ (:���S.�S as��������'9KX&L�EXE��9�+�!1�-eR,MPHASOE  k%�#�R�]!SHIFTME�NU 1:�+
 �<\�6//���� �!/Z/1/C/�/g/y/ �/�/�/�/?�/�/D?�?-?z?Q?	LIVE/SNAPn3vsfliv���?^3�� SETyU�0�2menu�?��?d?)O;OB��;����	(H'O�Oh\����� ��@⹭A�B8`�`��������A�B��C���G ��KSFME��0����� �M�O�<��z��W�AITDINEN�D���Q@WOK C �X[]��w_S�_�^YTIM�����\GH_�]j_�[�_�Z�_�Z�_\XRELE��gU@T����AS_ACT�0
h�a:\X_�� =��b�%  OLGE1�25.	r000y1��bRDIS�0��oAPV_AXSR&G`2>bJ<��O���Gp4 _IR   ��᥀������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� ��2�D�V�h�z�����Z7ABC31?bI�� ,�=�2��ܬ¯������
��Y���M�PCF_G 1@S}0A�������ҿ��`����,�b�MP��=AbI  �@��q�:��Q8|O`����t��Ϙ�?�T� ������D����k�-��߰��ѿp������� ����	�l�E��i�{� �ߟ�R�\�n߀ߚ�� ����2���e�w��� ��������.��d� =OZ�s�@��\ �����'9�� ��Tf����� &�/5/�\/ /�/B/T/f/x/�/�/ F��(?:?L?v>���u�(PBS{j�P_C�YLINDER �2CS{ ��&? ,(  *�?�=��#�?O�?8OM  �/nO�O�N�?�O$O�O �O�O_RO3_E_W_�O {__�O�_�_�_�_*_0oof�R�2DSw�a �"�hoxl�s�/��o�o�o��o�o�1�qA��o*yo�o` �o��o}�	�� ?y&�uJ��Z��� �m����?��׏��_�4�F����2SPH�ERE 2E�=� o_���_��͟����_ L�'�9�i_]���⟓� z���������F�X� 5���Y�@�R���֯���ſ׿N�ZZ  �$��4