��   �P�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�RYRUN_T   � $'�ENB 4 NU�M_PORTA �ESU@$ST�ATE P TC�OL_��PMPM�CmGRP_MA�SKZE� OTI�ONNLOG_IgNFONiAVc�FLTR_EMP�TYd $PRO�D__ L �ESTOP_DSBLA�POW_RECO�VAOPR�SA�W_� G %�$INIT	RE�SUME_TYP�EN`&J_ � 4 $($FST_IDX��P_ICI0�MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI�  xMKR�-  $L{INc   �o_SIZc8x�� k. , $USE_FL�4 ��&i*SIAMA�Q#QB6'oSCAN�AXS+�INS*I��_COUNrRO��_!_TMR_VA�g�h>�i ) �'` ��R��!n�+WAR�$}iH�!{#NPCH���$$CLAS�S  ���401��5��5�6/ �055������c����\1l5�1071p5��%VA�G���<�0TP��?��A5I2.L;c ��"��	AU$��Y4d��Y34	A[2)Y3�Y4-D� &H��&GH\0pAhF	~ChF�CRhFÞChF�n@�fH�̾ChF�n@�fH��n@�&GAA4B�D!Bz08�H`0Q�Fhz0�i�Hl.S�Fyz0���H�z0��H�z0�j�H�z0�&G~SxV~P�HU@�QxVVa@2vX9~P;vXUA~PPvXa~PxvX���SxV�~P�vX��cxV�~P�vX�@%�vX�>cxV�~P�@RxV�^c(E\0P,hf=@+fhC�chf�H# �5maL�chfQ�# qfhAP{fh�D�chf�# QPhf��c�hfaPqPhf�@�2fh�# Eh�>s(Ea�@PqHvP3Fx�7nsHv�0�qHv�P%sFxw�sHv��sHvf!`�Fx1p�&G��@�q�v �s�v1��p�P�vV�p�P�vvR�p���=AD��G&�aM���U=AAP z&��^�)�����&���~�)��q�&����
&����&�ae=A����eU=A�A�&��X��@(� ��@P����P ���J.�����P@����PP���`H U��en���u ��U��U������ �F&�
n@�P(���DB���z0��?���`�����6W?05�V1 �FOLGE���U�U  0h�M�AKROa�SU�CH�eh�BIN����D�o { �2L; 4%F|�SP��ׯ��J�ZDƦ�U
�  </t�̠eu>��  h=eq%�H��3Ʀ4A���5-��Y�}1Ʀ;2����="k���6��⯐�<uu�  amu���UB����"����tL?�������P$��"�X �01\0��0tt* _��q��F������ �,�>�P�b�t߆ߘߐ��m9}1��s����B�qBqu)w H��Iqs��{Zr��\tt���tt}1�'�9� K�]�o������p����7� 2t� ����� &�8�J�\�n������� ��������i7�, >Pbt���� �����(:L ^p������ � /$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ //2?D?V?h?z?�? �?�?�?�?�?�?
O? .O@OROdOvO�O�O�O �O�O�O�O__#O<_ N_`_r_�_�_�_�_�_ �_�_oo_1_Jo\o no�o�o�o�o�o�o�o �o"-oFXj| �������� �0�;T�f�x����� ����ҏ�����,� 7�I�b�t��������� Ο�����(�:�E� ^�p���������ʯܯ � ��$�6�H�S�l� ~�������ƿؿ��� � �2�D�O�a�zό� �ϰ���������
�� .�@�R�]�v߈ߚ߬� ����������*�<� N�`�k߄������ ������&�8�J�\� g�y������������ ��"4FXju� ������� 0BTfx�� �����//,/ >/P/b/t/��/�/ �/�/�/??(?:?L? ^?p?�?�/�?�?�?�? �? OO$O6OHOZOlO ~O�O�?�O�O�O�O�O _ _2_D_V_h_z_�_ �O�O�_�_�_�_
oo .o@oRodovo�o�o�_ �o�o�o�o*< N`r����o� ����&�8�J�\� n���������ڏ� ���"�4�F�X�j�|� ��������֟���� �0�B�T�f�x����� ����˟�����,� >�P�b�t��������� ǯٯ���(�:�L� ^�pςϔϦϸ���ջ� ds
 �q����t ���"�4�F�X�j�|� �ߠ߲�����ٿ��� �0�B�T�f�x��� ������������,� >�P�b�t��������� ������(:L ^p������ ���$6HZl ~�������  /2/D/V/h/z/�/ �/�/�/�/�/�//? .?@?R?d?v?�?�?�? �?�?�?�?O?*O<O NO`OrO�O�O�O�O�O �O�O_OO8_J_\_ n_�_�_�_�_�_�_�_ �_o_4oFoXojo|o �o�o�o�o�o�o�o )oBTfx�� �������% 7P�b�t��������� Ώ�����(�3�L� ^�p���������ʟܟ � ��$�6�A�Z�l� ~�������Ưد��� � �2�=�O�h�z��� ����¿Կ���
�� .�@�K�d�vψϚϬ� ����������*�<� N�Y�r߄ߖߨߺ��� ������&�8�J�U� g߀���������� ���"�4�F�X�c�|� �������������� 0BTfq��� �����, >Pbm��� ���//(/:/L/ ^/p/{�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�/�?�?�?�?�?�? O O2ODOVOhOzO�? �?�O�O�O�O�O
__ ._@_R_d_v_�_�O�_ �_�_�_�_oo*o<o No`oro�o�o�_�o�o �o�o&8J\ n���o�o��� ��"�4�F�X�j�|� �����ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ǟ����(�:�L� ^�p���������ïܿ � ��$�6�H�Z�l� ~ϐϢϴ���ѿ���� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r����������� ����&8J\ n�������� ��"4FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�//?,? >?P?b?t?�?�?�?�? �?�?�?�/?(O:OLO ^OpO�O�O�O�O�O�O �O _O$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o_2oDoVohozo�o �o�o�o�o�o�o
o 'o@Rdv��� ������#<� N�`�r���������̏ ޏ����&�1�J�\� n���������ȟڟ� ���"�-�?�X�j�|� ������į֯���� �0�;�T�f�x����� ����ҿ�����,� >�I�b�tφϘϪϼ� ��������(�:�E� W�p߂ߔߦ߸����� �� ��$�6�H�S�l� ~������������ � �2�D�V�a�z��� ������������
 .@R]�o���� ����*< N`k����� ��//&/8/J/\/ n/y�/�/�/�/�/�/ �/?"?4?F?X?j?u/ �/�?�?�?�?�?�?O O0OBOTOfOxO�?�O �O�O�O�O�O__,_ >_P_b_t_�_�O�_�_ �_�_�_oo(o:oLo ^opo�o�_�_�o�o�o �o $6HZl ~��o����� � �2�D�V�h�z��� ���ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n�����������ڿ� ���"�4�F�X�j�|� �ϠϲϽ�Ͽ����� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p���������������� _ds
o�qu���q����qss���^�tr t��� q �t ��CUgy����������`��J� L K Mq�uqs)A�rskq)o �t!'�tt1K]o����������akds���,�rK8tB,  u(�H""I Z  \9J/\/n/�/�/�/ �/�/�/�/��?"?4? F?X?j?|?�?�?�?�? �?�?�??O0OBOTO fOxO�O�O�O�O�O�O �OO_,_>_P_b_t_ �_�_�_�_�_�_�_o _(o:oLo^opo�o�o �o�o�o�o�o o 6HZl~��� �����2�D� V�h�z�������ԏ ���
��'�@�R�d� v���������П��� ��*�5�N�`�r��� ������̯ޯ��� &�1�J�\�n������� ��ȿڿ����"�4� ?�X�j�|ώϠϲ��� ��������0�B�M� f�xߊߜ߮������� ����,�>�I�b�t� ������������ �(�:�L�W�p����� ���������� $ 6HZe�~��� ���� 2D Vaz����� ��
//./@/R/d/ o�/�/�/�/�/�/�/ ??*?<?N?`?r?}/ �?�?�?�?�?�?OO &O8OJO\OnOy?�O�O �O�O�O�O�O_"_4_ F_X_j_|_�O�_�_�_ �_�_�_oo0oBoTo foxo�o�_�o�o�o�o �o,>Pbt ��o������ �(�:�L�^�p����� ���ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ�ſ������ &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt �������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�? ?2?D? V?h?z?�?�?�?�?�? �?�/
OO.O@OROdO vO�O�O�O�O�O�O�O �?_*_<_N_`_r_�_ �_�_�_�_�_�_o_ &o8oJo\ono�o�o�o �o�o�o�o�o	o"4 FXj|���� ����0�B�T� f�x���������ҏ� ����%�>�P�b�t� ��������Ο���� �!�:�L�^�p����� ����ʯܯ� ��$� /�H�Z�l�~������� ƿؿ���� �2�=� V�h�zόϞϰ����� ����
��.�9�R�d� v߈ߚ߬߾������� ��*�<�G�`�r�� ������������ &�8�J�U�n������� ����������"4 FQ�j|���� ���0BT _x������ �//,/>/P/b/m �/�/�/�/�/�/�/? ?(?:?L?^?i/�?�? �?�?�?�?�? OO$O 6OHOZOlOw?�O�O�O �O�O�O�O_ _2_D_ V_h_z_�O�_�_�_�_ �_�_
oo.o@oRodo vo�_�o�o�o�o�o�o *<N`r� �o������� &�8�J�\�n������ ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϱ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������� &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/��/??0?B?T? f?x?�?�?�?�?�?�? �/OO,O>OPObOtO �O�O�O�O�O�O�O�? _(_:_L_^_p_�_�_ �_�_�_�_�_�Oo$o 6oHoZolo~o�o�o�o �o�o�o�oo 2D Vhz����� ��
�.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� �8�J�\�n������� ��ȯگ����"�-� F�X�j�|�������Ŀ ֿ�����)�B�T� f�xϊϜϮ������� ����,�7�P�b�t� �ߘߪ߼�������� �(�:�E�^�p��� ��������� ��$� 6�A�Z�l�~������� �������� 2D O�hz����� ��
.@R] v������� //*/</N/Yr/�/ �/�/�/�/�/�/?? &?8?J?\?g/�?�?�? �?�?�?�?�?O"O4O FOXOjOu?�O�O�O�O �O�O�O__0_B_T_ f_qO�_�_�_�_�_�_ �_oo,o>oPoboto _�o�o�o�o�o�o (:L^p��o ����� ��$� 6�H�Z�l�~������ Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲߽� ��������0�B�T� f�x��������� ����,�>�P�b�t� �������������� (:L^p�� ������ $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ ��/
??.?@?R?d? v?�?�?�?�?�?�?�/ OO*O<ONO`OrO�O �O�O�O�O�O�?__ &_8_J_\_n_�_�_�_ �_�_�_�_�Oo"o4o FoXojo|o�o�o�o�o �o�o�oo0BT fx������ ��,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��� 6�H�Z�l�~������� Ưد�����2�D� V�h�z�������¿Կ ���
��'�@�R�d� vψϚϬϾ���������*� 