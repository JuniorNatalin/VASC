��  	��A��*SYST�EM*��V8.2�306 4/2�
 014 A�5  ����A�AVM_WRK_�T  � �$EXPOSUR�E  $CAMCLBDAT@ �$PS_TR�GVT��$X� aHZgDIUSfWgPgRg�LENS_CEN�T_X�YgyO�Rf   $C�MP_GC_�U�TNUMAPRE_MAST_C�� 	�GRV_}M{$NEW���	STAT_R�UNARES_E=R�VTCP6� %aTC32:dXSM�&&�#�END!ORGBK!SM��3!�UPD��ABS�; � P/   $PARA� �   ���ALRM_REC�OV�  � A�LM"ENB���&ON&! MDG�/ 0 $DEBUG1AI"d�R$3AO� TYPsE �9!_IF�� D $ENwABL@$L�T P d�#U�%Kx!;MA�$LI"��
F �APCOU�PLED� $�!PP_PROC�ES0s!�(1s! �(�!> Q� �� $SOFT��T_ID�"TO�TAL_EQs �$0'0NO*2U SPI_INDE]�?5X�"SCREE�N_NAMr ^�"SIGNe0�/|�+!0PK_FI� �	$THKYޛ7PANE24 ~� DUMMY1d��4d!�54�1���ARG�R�� � $TIT�!$I��N D@dDd D�0D5�6U6�67�68�69�70�7G�1EG�1E�0G1:G1DG1NG1�XG2cB�1SBN_�CF>" 8F CNV_J� ; �"L �A_CMNT�?$FLAGS]��CHEC�8 � E�LLSETUP �	 P� HOM�E_IOz0� %�5SMACROARR'EPRJX{0D+>0�dR{lTD�AUTOBACKU��
 �)DE7VIC�3TIc0�A� 0�#��PBS�$INTERVA�LO#ISP_UN9I��P_DO�V7��YFR_F\0AI�Nz1��1�S�C�_WA�T�Q-jOF�F_� N�DELZhLOG�R�1ea�R�?�Qf`�3?��� {1�5� �MO<� ZcE D [�MZc���aREV��BIL�g���AXI� �bR 7 � OD7P�a�$NO�@M�t�cr��"w� u<q�x�`Z0D�C �d E RD_E��`Ts $FSS�Bn&$CHKBD�_SE�UAG G��0 $SLOCT_�V2�q� Vzd޾%���Q_E�DIm   ȫ cQG�CPS<:`a4%$EP1T1O$OP^02danp_OKnrUS�!P_C� �q�T�vU ^UPLACI4!TQ�?��p( �QCOMM� e0$D;�Q�J0�f`�y�?�2�B�L%0OU�r , K�QQ2QU B�@y �O]Å��CF�Wt X $G�R� ��MBZ`N�FLI���0UI�RE��$g"� SW�ITCH��AX_uN)PSs"CF_��G� � 
$WARNM"`#!�!́p�@LI�f�NS]T� COR-�R�FLTR`�TRA�T;PTb�� $A�CC�Q��N ��r�$ORI�o"�R]TlP_SFgB��HGz0I��bT��1�IʐT����K�� �x i#
Qnr�H�DR�2J; �3I�2�D�3D� F�5D�6�D�7D�8D�9�"���CO�D <�F �����#�܀O�_M�� t� 	PEq0�1NG�1iBA� Q���q ��!�Qp�0=q�0�I�P�PJ���G�S��pm �RC ��4���"J��_R��g�C��J����ļJVep�%C�X���p0�h ��AzOF�� 0  @F RO0��&9�6�IT3c9��NOM_yV�lS� $��D Ԁ0��A�B�'&�EX��B0��P����
$TF�E0��DM3N�TO�S3U8P�+� -0P_H��j 1�E{� �%�Y#&�d%(��1d�$�DBGDE}!m_p$��PU��1a2)��I"���AX�Ae$]eTAIn�SBUFivY�>/ � k�f�[PI�$��P��EM��M��^���F���SIMQ� �$wKEE:�PAT0������N#��Y"�$�L_64FIX/��L⥟TC_��� ����c��CI됎�PC9HOP��ADD��� ������I"m0p�3�_��!f���n!
�`�a��W���d"�$��MC�� �0yJBE�ͤz��l�+�i�s ��� ��p�CH� EMP�#$G�����p_�lS��1_FPm��@��SPE��lPn�������� V�q<r�A̛�JR�<rSE�GFRA��3 �R>�0T_LIN{sM�PVFs!#�'�_��"�#m�"� R��|$�y� D )�� �`�����2�f�)P����Ţq�f�SI!Zc��T����3�RSINF ��G�R �e3 e��> L�з�gCRC(�AcCCn���3 ���*���1M�a������D�&�e#
)C+e`TA�M ^�&�T(EVTT&i�Fj!_F���N�&�@f�`�((��r����'�\j91���A! �>p��F-�RGB�ª�FB �ׂ��De�R��LE	Wر�Q����/��.  ���Xs"� ��Ư�5b��#�R� HANC�$LG~��!�QU�y�gp��6�A:`� a�c�R?2 �3p0��3�\��8RAnS�3AZ���7HP ��O�FCTC�Y07�F)����\R�ADI�KO�H @�@�o��D~�.���6�S�p����qM�PW*���M�4A�ES��l#���0I}_�4#  �=I+$�CSX��H�B��$*�?p�s��T�B��C�0N�p�IMG_HEIGHmq�rSWIDK��VTt��M��pF_A 8{��B`EXP�A4�N�U�CU7�]�U%�w% $_�TIT���r�s�p��E�:RZ_% {�&*�b{� ��A~�NOwPAD	q?W�i?�,������DBPXW�O�&�'��$S�K���r  <�`T�0TRL%�( ��,�A!���@��rD�J��LAY_CA�L�q	��`�@�gPL�	�G�SERVED W�wb�w��'��T	���9��0����`dAA%�)�b��PR�? 
8�D"����%�* _���$��$"L�L2oy+|"ѐ��&�y,�"��PC%��-�p��PENEL���!.�"�(OqsRE}��r/H�0�C�� *$L2�+$os��+@C�T 4��O�0_D�A��RO����䤍�>|�RIGGE��PAUS��VET�URN���MR_��TU>��a�E�WMF��GNAL����$LA-��n��,$P��-$P\@!�.�b��1C!�!��DO` ���\�H��b�GO_A7WAY8�MOD�0~�B�DCSrp�EVIm� 0 oP $іRB��
�PI���SPO��I_BYT2�����TXw�L$�1 H�� 7��Ф�TOFB��FEl������lw�CU2�DO����0MC��N���7�(`����Hy@W����w w�ELEGR�3 T����cCINQKh�����U�L��cHA��}$��} w�����w4 ��`MDL��O 23��(�O��^����C�2����J]�}O�m�}2�U� r�h�������	������%U5� $ ]��0�PcC�PZ��Pa5�бw��ϲ��̵I!DJ�˶�b˶W ���gNTV��вVE�Ր(РW�D�2W��J�&���pSAFE�)���_SV�BEX�CLU�a��>2ONL���Y6��3x@��Qw�I_V�@�PPLY_���� Ƕ���_M�"��VR'FY_�c��MS3�P!O��x@!֧@1~S4ӂ^�O���İ��@� 36��`TA_ ���  v�_�SG�  7 ��CURπ�}S��8tpUQO�REV�ٯ���jPUN�p��ԥ��Ё�����0���Ѱ�@����EFаI.�r8 @� F���T�OT�At<�At�'qAt^� �+�M���NI�r9 L !�`��Aʱ���DAY	�LOADИ�6tv�Bs5>q���EF�P$�X�:�d' SO����\��`�_RTRQX�; �D�!O��RQ{ ������:| C7 񙔈�A;`���< 0�Z��p�Z�L>��6DU5��b;CA�� =9�[`�NSk���ID� P�W93U����V��V�_U��< �D�IAGr�u>8O *$V��T%@ep
p}R�rt��{V2`��SWB��u���R �2�;�� �OH�r�3PP2a}IR�Q}B���m������	��BA����D@�H�����=��CY ގRQDW�MS�� AZ`w0{LIFE�`�/Hq��NB�K��@��!�����C�@f�NrЀY0�QFLA�4��OV�@W.`���SUPPO�`�Aĝ��`_���z_XP�C�a��Z�W���A��B���CT�%U? `��CACHE�'C"ۣ�կ����� SUFFI��ϰ�`%a6t��Bs6�>q ��DMS�W%U@ 8��KE�YIMAG��TM�F�C�!с�&INP�U}R ,�G�VsIEL �1A ��BGL/đ��?�� 	dnpfPcB0MP�!g1IN^�Tb4��	UBv�JB�a�dJ��O#QT�3��S��Uu59d�;��OFz��H��C �Va!gOTF��ץ1�D>[�P_GAI�Q��p�@�@̒��NI_�0�C���5���6�PTIC��O�PE���"���}1�A{�PCF�@IN�y��P[EAq�@!� ��A$P�3D�  P��6D�7I��8T�=�Rv�=�AVE�FFBP�c�C���3AW_�@<��E����DO<4S�LO���1TERCE/���DL/`�J3UFU'RQ�E�e{0�Px�E}1�DX�B�FE��3N��3qPQ;`��5�R�6�R�5t��G�FF� 䠣�$s�2��G �1�0���1F����0�3��0 ��AbB��cCGARRg#i0�9T$ 0<2%cyftqRD_4�0&6FSN�p��T� �F�SY��DI"e�CH��A�D��dEG<�R�F 	h2u0��Hb�C9�0ǰY����1�@3�G 9�2A I� {  _��3]6�0�s�1�s�1��r��D Ц$J��z�STp@! �r)��tk��tv��t���pEMAI���/1s��� �@AUL��qK�")8}1COUdP䙀-!T!���L,ȍ@�M�SU��IT h�RZ�U'}�N��F 'SUBRT��C봅�8�*rw�SAV~�@� ES��m�������9P��M�ORDM�p�_RPd���ډOTT���A��P�60��s�F�AX��,��XRP��TDYN_�>�M�b��6�௕�G3��@IF� �����b=�N� �05��r�C_RO�IK�"���Ҟ��@�R�!���8��DSP$�&��PA��I(v��H�ß���U���D���M�pIP0Á��D�  ڔTHRES��`˕��TZۓHS@�bۓR`�E[@��V�����@�㑤P��NV���G����]�ؖRPF�B��d���@(��!S�CbRu��M-P��F�BCMP�À�ET��a��O�"FU�D1U'��QPPEP����CDљ[���-3h�~� NOAUTO��P�$z���z���PSy�CR���C<�BE &�v����QH��в��r� г���@N����S�� k���v��������!��7��8��9��B����1�1�1*�1�7�1D�1Q�1^�1Jk�2y�2��2�U2*�27�2D�2Q�U2^�2k�3y�3ʩ3��3*�37�3�D�3Q�3^�3k�4�y� �v�OUT|� ��R � "@�	WvPRuPLCWA!R+v�`����R��$FACm�SE���$PARM1��2m�"k��$x³�pA�P$�XT��!S <�)9I�g�0Rv���枵}@FDR~dTT @  ����E-�BE�11N(OVM�4T�A\�oTROV\�DT��|�MX��vP&�{�N��IND��:
���`E�PG3���� pb1�`DRI�@�c�GEAR�1I%OQ�KL��N�@:EFF\�k�� �M�Z_MCM1�E<��F�UR5�U y,��V�? �F0@?� Ð0�yEi@� 	(�p���2� V�RTP��$VARI�5TD����UP2_ 3W *�?�TDI�iA�>�TV��  +�H�BACG�X �T�p@�U�=0)$/PROGC%?���:�b�IFI�� �wYPa��!,��FMR2�Y ,�k��B-�Mp� 1�8J\s�}0p�L��_���AC@IT_<[U�C_LM��>(DGCLF����DYt(LD���5�������
đ�uZ�� ) T�F9S؀�t[ P�P�"|:2�$EX_�!��(�!1'�נ���!3�;56�G���\� ���2��4l�ON�����1�T�1Q�GRt��U��BKU��O1�� ��P�O��9�0$�W5�0M�6`LOO��1SMzw`E�� �����`_E ] \���  �,PM�5�^�9ORIp�1_>�7�SM_M	��0`�5�)P�T�A/Ia!IUP:P ?b� -��b�]$�5v@^��G�{J� ELTO�CU}S�@ONFIG����A� c1aCrD_$9U+aא$}��A��@P� OT�G��TqAk�-�3SNSTv`�PAT`�f`RPTHJ(�N�E� ��W��BARTE`�E�p����r�AR[pRY��SH�FTR��AQCX_SGHOR1�K�.F 9@�$HG�Pa>!.�OV�R����PItP;$Uz�� M�AYLO0� !A��`� ��Q]���]�ERV��Q���Z ���Gv`QR��t;e���tRC���ASY1Mt����AWJ�G����E�?QkibQ�U��d@A�CU�qP�YUP���Pġ�VOR@MF��?0�1 �c�r��2�6P�@!P����q�%d Ƚ�x.LTOC�A�1i$OPo"���(�2��pH�O��Z�REbpRأ��)�K�ReipRU�u}x|[QDe$PWR$ 3IM�ubR_Xs8TgVIS/@�bT,r��B e� $HzC!�ADDR��H�1GR/�$����v�R3�����f H��S��N���\���\���\�*Â�N�U���HS[�MN�!g uB�trq�[�OL1��h���<^��0ACRO�p�AhqND_C1�|�a<�tšROUP��!rE_ÐI1�Uq"q1�� 6�2��<���<�Q�=���<�*�<�7�6�AC&��IO��D7����G���� �h $� Pp_D��0�⣂�PRM_+��H�TTP_|�H#�i{ (��OBJE�l��t$�LES(����ְjN0����AB_��T�3P�S|����DBGLV1��$KRL�yHIT�COU@�1Gf�L�OC�O�TEMP�t�����zpv{pSS����HWe��A#��kW��`INCPU���pIO�e����r�����*�,�oIBGN�$l����� WAI�s�aP0����R���FW$ ېLOm��s|���vy�AN�A$Bo��������������RT�N/`�CUF_DA�TA�㖠����_M�G�2/ F�>�S(SE8��r��8REC���MN�b�2�h�I� m @� N�_�h�Y�3t���EXE�wɒ�Ф _�X�u�0�n�$SC�H�`�QP�R��F�LGvQ: 2�	/�o`o�����v ��OP�8��1~�TRA�B���CS8��9�p�x $C�CTA���'�IGN�M"oO҈0�M~�T�����v���vN_PC�SO�QUp��ECF Ba��Q���u��Ғ�	�\r��L�������@D�FRs������SPTx �$���SEQ_� Z3NS��H�*�ɀ��rC�q�@Xl�S L�}Pr�Q �-@o�bc���0�se:!X�IwOLN4q 8��R�$SL�$INPUT_��$�p��P- ���&��SL���!rr���#����ݐF_AuS�"s:$LO $�O��Р�r+������PHYP���^� �8�UOR��#t `J��(�%�s�%�|���pP�s������|������ ���UJ}R�u � 9N��UJOG�G${DI,�$J7�VdJ8O	760I�A|Xj7_LABQ�HpZ �NAPHI�� QY�D� J�7J8�0_KE}Y� �K)�ML�%v  �AVއ�P�CTReS�F�LAG:2��LG�$w �����~Y3LG_SIZJ���0>� =A�=FDHI<S�1J;@ =:tsC�� �A��j�@�X_R��������5��LNCH2x����U01#��!BpU�)!(��L2#("DAUN%E�A�)�Dtd"Z GH�Er ��M�BO}OQ�yt Bd��pIT�Ø${�e�#�N�(SCR��`�D��|[2$�MARGI�D�,�X�ct2��M�	S0�L�W�$M�=$X��JGMC7MNCHL�M�FN�F6Kl7q�j9UFx8�Px8n�vx8HL�9STPx:�Vx8àx8� x8RS"�9H�`�;U�C�T�3 �bX�p7CIU䑌4@7�R,6� +�2G\9lPPO�G�:�%�3Ԇd2OCG�{8���GU%Ij5I�3�B(3 S43Sh0l1�P�rC�9��&�P�!N݁-�A�NAM�Qq�QVAI|� �CLEARfDn�HId�~Sr�~R5O�XO�WSI�W�XS�X8lҸ�i�i1���Tքn�DEV��}�!_BUFFq�z� �pT0R$�IEM����' Q
bjqq{� �pp���ˁIpOS1je52je3ja 	c~Q	p| �! ߈�aZSq��{���IDXtAP�ƞ@z�jK�T���Re Y���a {$EvC{T�㐜v)v ��ch�} L�s������`�����w3��u�Kc~�#_ ~ �� +�#��!�s��M�C" �! C�LDP��vUTRQLI� wT2 �y�t�� ���p͑�nQD���ڠL���t�ORG2 B!�'���������!���s͔� �����tE�t�SV�_PT�p��R�Ǆ>φRCLMC݄m����]\�MI;SC� d%!�a�RQ����DSTB��` K��!X��AXvR� [�t�EX�CESm *4R-�M��⡂��?��vT 
X-��㠃
�M�_�I������r�����MK��c \�P�MBۢ�LICL�B� QU�IRE,CMO>�O�N�DEBU��
�G�ML���Ш���e�H�Pށ ԇ�2�Di $�D�$U�PyACKE�D����DPxv��IN�b$q�_Q �pI� U�������/�	��=�U�4�T�I�,�ND:!SSb�#""$f��DC�6$IN]ю3'RSMD ���PN�r�BC���y�P{ST��� 4q�;��fRIl �e�e�ANG�bI�P���AQ���;�$3ON,"�MFq T��i��00�uz� 3��SUP�� ��FX&�IGG�! � �ဃs��#�s6F�tR{�v��b������ȵ�����+�DAsTA���ETI8 f,��1�1`INb�� t?�MD?�I�n!)M���YӇ�U�H8#�SX�DIA�Y�ANSWe�Y�Pa�A*X�Dl#)Oŀn��� ��CUSqV���I�T���LOf �������G�0��5����� � ��RR22��O� ��J!Á� d$CALI�Q��GrQD�2f`RsIN�0G�<$RR��SW0�����AB�CS�D_J2SE�e�I�L�_J3��
���1SPm I�P�����3���ѓ�I�B��J����āOa�IM��CSKP �z<�- kS<�Jm!��Q<�m�S�m�c��_cAZ˂	��ELa<���OCMP&�����1�� ���`1����� ��Z��0�OINTEVpSb����2I�Vp_N²��7�a'�43̒�A	DI��(�`�DH��6 ���Y`$VQ঳�a$l1$ �!�`��Q�-�2��H �$BE��|�	�qACCEL������ IRC_9R-��ONT�a�c�$PS���rL  �!�s -!sPPATH�	Z�"Z3)����_ga����ʂ�C��� _{MG�Q$DD�<�"$FW5�1�`�����DE��PPABN1ROTSPEE�ka/8�pc�kaDEFۑ�~)$USE_P�J>SP�C�@>SY
 �� ʁ �aYN1�A�c�x&,�o�x!MOUf�NGtB�OLJ�$INC�� ����X��'3�Y�ENCS�P��I�!�V�IN�bI)52�΃c��VE� H�*223_�U>��<3LOWL��Qz@���p�%\6D�]@I�3� �p�%�C�' #6MOS�P�M�O���`ʇPERC7H  y3OVp t" �7�a�3��_2̈́���� ��b%��P*�A)EL=T*��)�$5��_:�ZFu6TRK�4�bAY��Cܑ�A)�E�C8!��`�RTI���"�`MOM�BX�ܒc���G��D��C\jb� DU2��S_BCKLSH_C) U� �6�0�#��:T�"xEZ�!e�CLAL2`�"2���@�`wUCHKt�p�eS� RTY��B�5$�U�0�_�cN�4_UM���YC�SήSCL�T# LMT��_Lg����T�gE m!`k�Pe���0Q�!&@bd�8P	C�1�8H�pl���U�C뀎rXT� �C�N__�N���f�S	F��9Vb""�7�p�a)u�hCAT�^SHo�_���&U�Q�6��*����PAL�T�"_P�U�C_�p��P�F�0�q�C�t�UJaG�����sJ0OG�g>�BTORQUT �� �3�I�/��2�A��_W�E�D��7���6��6�I>�IL�I�F9�)��#��VC� 0R�䒬�1ಎ��Əc���JRK������DBL_�SM�!5BM��_D9L�5BGRV=�6�0�6���H_���]d�COSq��@q�LN��������� ��� ��h�Қ�����Z���6�MY���}��TH��1�THET=0e5NK23�[�l���CB`�CB�CT�ASƱ��h������`�SB���k�'GTSE�#!C�� ����|s���ϓ$DU�P>G�D��!����3��AQ��&�$NE�B��I��#���L$~ O�AS�|���c�n�n�LPHq�Z�45Z�S��ͳ��ͳϕZ�ޖP�����~ V��V��T� ��VźVһV�UV�V��V
�V�H�����µ�:q��һUH�H�H��H
�UH�O��O��OI٪��OźOһO�O��O��O
�O��F�Z��������ԑ�SPBALANCE��~aLEȠH_S�S�P��4���4�ϖPFULC8�_�G�_��ϕ!
1���UTOy_�P�uT1T2���2N�Quc���O@�Aa�?�0��ATK@�O���'�INSE9Gu~1REVB�~0�1DIFtEF	1�l+�r1�g@OB!�gQ@��G2����Q�?LCHWAR
"g"�AB�q�E$ME�CH�� ��!��VAX�APEd��u������ 
����5ROB�0CR)���b� W��MSK_|��� P ��_R R���+:!vD1r/0-"+ ,3ET+ ��IN��MT�COM_C��� ��  �3� !�$NORE3���OPWO��� �w, k SBU఍�QOP� �T��
U�=PRUN,q�PAR D���\��0_OU�!��S�AB�"$ I�MAGVQ( B�Pf�IM� BIN'��BRGOVRD<��	@P!Ap�!_��q��R�`R�B�`��[aMC_�EDT_� K`N�l�M�JaPMY1�9IaH�nSL�6�" � x $�OVSL��SDI0DEX�c&�cKA "V�!$N'!��5 %#:'5(�p��_� �" � @@�pl"���2� SB
&�_���'�!�! ���0�ECT�  ǚ H(��PAT+USP{@CD�Z;DX�&BTM�'�!	I	�4Ia�#�" � D( E"�"�Z�E4��!FILE8J@gP�!EXE� �Q �72K24t#�{ ) �� UPDATZ1$T�HXNDP���x���90�PG7��UB�!����!�!�#JMPWAeI'pP*#�5LO`¤F�p�!�RCVFAIL_C�A��1R�@� �V�a�dx��<E�R_PL�#�DBTB�q�UBW�D.F� U�P/EIGpI��TNL#p�0D�BRT�� ERcVE�c�D�b��1�DEFSP�P � L( ���@``�qp�CUNI"7�@b�1RR0!�.�_L��P�! ��Pr !� 0�q�!N] ATA$�uNP�gKET$R#�BUt�PIPB!� h~�ARSIZEp�@E0GQ�RS� OR~�#FORMAT���uDCO�Q�EM2���TSUX� :" ��PLIpB~!�  $| �P_SWIp�%�����U@p@AL__ � $�AAV�B���CVD	�$EZ1�`C_�zA� � � 1Q�VaJ3��V�80RTIA4hi5�hi6VMOMEN�Ttc�c�c�c�c| B @ADtc�f�c�f�cPU��NR�d�e�c��e�b �T�?P H$PIQ�� 6�H�Z�l�~���!ڦ������� ��GQ�&S/PEED�G�R�t E�D�v�DE�,@�v���x��y�ESA�M#��F��wL�EM?OV_AXI�!��z��%���7�z��@1d��2dR	 md��0	`a Б�INڌ	` /����؄B�#���<#�C�GAMM��A�܋R��GET�rFI�MS�PDcd
��LI�BR�1�BI�@bS$HI�0_^� f��E`ŘA���ӖLW�� ����$�Ӗ?b���@aCfEq�|��  $PD#CK����_.��PdւSiaɅ���c����f��c �+$I� R��DW���1"D��LEa�q�!��?hᠣVpMSW�FL1DM`SCR�86�37��U��q� 	+Pq]�p��P��URB���G�R��S_SAV�E_D����3NOC`C�!�2Dd����Sj <v幾Uy�mp���@�pW�v<Ƚ�.aO�AA��񊅰���e�x ��vv��ǜ�ZÌ���1 ��QMu�o � ��YL5s ~�ɇ��~�����NB�KA���WѰ�(Ղ�4��`�����M���L�CLK�aD��^�1j�8�PM��� � � $����$W�Є�NG1]a��d��#d�� *d��1dV@��s���S���	`XPO+caZp&��P@t� p�| ��Uv������,�;�Ca_�� | �Si���i��c��c ��mj	���jE@��� 
���y�� t^`��P�Q�PM4 �QUP� � 8�8PQ�𽡤QTH� HO��HYSf�PES����UEr����hP��� � �6B;Q#��#��_`� 'Ѵt���EN/	PBG_@B�[mB�?�#*#Jہ��I̢�pEW �vGTqF-b"�PO�4�   �𮗫"sUN� N� I�9O�rp� PD��E��-3�BROGR	A�!��264M ���ITh@�{ INFO�� � ������� =(àSLEQ�v6H�u6�x{ �D�0p�����Ov����#5��E��NU���AUT���COPAY���0��qʰM��qN��^�PRU����� gQRGADJ�v!�wRX'��B$PP&3�&W(P(`��$�s	 �3EXF@�YC���!N�S�T� �4AL�GOk�.`NYQ_FREQ��U �w�!�T�LAhC�!��b.��5CRE�0��l��IFQq�NAT��%�$_GhCSTAT�@4��M@R����31	���Q31��|$E;LE�0 �Nb�SEASIr1��� "�a2�1���6BƀI�a�"�q��M���2AIB�Q/`E� �pVU1�6BAS9b�5����qU�@� ��$�1�F$|$��� X� �2 2� 	����QFBPGQ$|р�eE|F z&P�Fe1�=GRIDd��SB|P�wTYs3;�| OTO �1Q)�m�� _4!E �B�wRO$��$� �v��LI:�PORAS��C'v�BSRV0)lTVDI�PT_�p@6PHT��RW�pRW4PYU5PY6PY7PY84Q���PFs�e1�~� $VALU�3����4��L�Q�$�| n5	��C1
1���0AN���R�1Rp�!��TOTcALQ���7cPW�#�I�AMdREGENKj`b4�X!G�s�&��fm�TRC�rKa_!S���g``�3V'����c>�1E:3�@��¸��cV_H�@DqA}��`pS_YƱ��&Se�AR}�2��>@CONFIG�_SE��`RJ5_ě �������D� �4{�O�v�k�F�P�S��F�f�C�_F��m���L�����(cMϰ���q��r^⃁z��DE�հ2�KEEP_H/NADD�q!��0�CO�0+��A�r%�,�Of�
���q�p,�1��,�REMC��+����Bh����U�4e+�HPWD � q��SBMs! �uB� ,àcFL�з���YN�p
�M:�C���pQ�Ern�� �l0DB�oMTRI�DA,��B� 0�K�TCLA�����U AYNS9P��֡SEAꠁҖG_P�Tn���Bο�RGIn�QSOCLUK ��P��L)a�$SC`0D�#ےALI�r���S��B#U�A}������� ���w1��_�P�H�TIC�[�`�p[�RE3VIo��OLP����p�FK��_F�SS#EGQ���b�,@�Tc3� �l0CP���TU� MSEC��MN���̢���H��`�0�G����0O��1�$N�̡_�e�$�PA� j�P�vO�iP��MLr P�� ~� ց|е��e1��  $OW-����G����p@���Hp2C�ĹAü(�!ߤX�AX�Q��A7HI��6���ٔ�2��Ϛ���B�V�EP���P �`Q���H�ߢ�r��V�t��`a�B^"�$4:�Q������p�MĢ�y�O��l""�SM�H��<�M=�2�� T�L`UP_�DLY��ÆDE#LAk�>a2Yߔ��� �QSKI�'�� �P��OF��NT\P�B��P�� ���`
��P���a�� v��l���vP�ڃP��@�P�ڝP�ڪP��9���J2#����yrEX@T�#z����z��.@�z���T��RDCa�� �s ��0TORq���	��!�����SD�RG��H��k���G�g��eER�qUBS�PC�G�z�?2T�H2N�!D�#�1�� ���@��11�� l�p2�F1�7��Ta��� O ѯ%��^�����SDx��VAHOME��W �]�2e��k��}��������� �
]�3e������\0B �]�4e��ew���� +�]�5e����p*< t]�6e��_q����� �]�7e����� //$/6/ `]�8e��Y/k/}/��/�/�/  ]�S�πf��  �AqX^�u`� (]�Z��ET�yp���m2.fk3IO�p�:I�0�� �]�PO}W�� � U0�K����]�(d s���2$DSа�IGNAL#gf�CxJ�2��S232q5'� ����%8��ICEt����³���ITq&aOPBI�T"cFLOWCpT�R003b��UXsCU:+�M�SUXTđ��I��FAC1Dų%@� 		@CHQԣ @{p�p��C�$�`�`OM,p_���sETޠ�sUPD�p]A3� �	@P�@��Q�� !�(�s�A�����)��.�EWRIOc��PT:p3T�2_���Q/PDAMV#WR���/9D��qV���6FRIEND(�@�UFi��t�P����UMYH�p@���G�TH_VTE�TI�R���R�P�XUFINV_���>��WAITI���W�X���Y7fG27WG�1��@1SQbbgpp_�RE�O_t��s�Q�`���[PC�C�u��_T�C3��Ķp�e<�G(ˀŲtqֱ@&Q/A��r�jQX�EV��Ea�������D�X s�ML����`@��SX��]E#T�CG3�IWCPgws�|tD�LOCKkuvӮ�V���q�ta�$�f[�֐�pkQe�qY1}XlP2*o[2�{3o[3}Z�y '�~Y�yC�6.�s.Цr$VV��V8eVDl�ь�a�b!�غ��F�sρ��fqB����`�R�ɠ��E�$߂�S�@a�Tu���CPR����uj�Sl�<G�� ��D�C� ����%s[��w���[���p�@|`�@���
p�DS�1� ؚ�R_6�oQ��7�o$RUN��AXSA��`A�PL�QV⮒T�Hb�J���6�aqT�F"�NT���IF_CHeS��~�qU��6��G1��0��Һ��6�_JF?�P�R�`���RTCw� ���GROf�&A�MBVq̐CrÃ�f�`UI#���BU)c�RSM}��a`r�_�W�P�TBC_P��PCM��D��ЖLDR��ރ�A��@��̮c�IT�"7���v��TA��� s�D��|� �ҙ��� ����� ݾ2�  2� �S��>g��	| �Vд��}�I�t�ˀ~�TO�T��~�D젖�JO�GLIzC
`E_P��qBO��}����`�F=K��_MIR��Ѵ2{`M>r�AP]q���E)P�ҔJ�SYS��˂J�PG'�BR�K�bѕߐ��I"1�  N�pSY�x�D8�A~��BSO�}���0N��DUMMY{15U�$SVVp�DE_OPoCSFSPD_OVRU��� LD��óOIR��� NP��Fߑl�Ʈ�OV��SF����.�F �́ճc�8ؿQ˂LCHDL>z�RECOV��[P���W�PM��vձ�R�OoC����_ И�s @�&`VER��_$OFS&`C;��SWD��r�����R,ū�TR�1W1FpE_FDOƃ�Ӡ��B��BL�����1K0%�V�A�B�@��b�2 �G�,�AM*Ã�0D�Z��t�_M0�|Bx��3��T$CA����DU���HBKX�AЖ��IOoU���1qPPA������������2��DVC_DB)c0�ё�21����́H�1P���H�3�P���ATIOˀ��A{���UtS젆6CAB��nR�c7p���`�S��A��_�@ЖSUOBCPU�2��Scp �0�B��@sj�B���2��$HW_C _ dЧs5�sAta����$UNITb�|\ U ATTRI��i��CYCLϳN�ECA����FLT?R_2_FI��8����6��Pǻ��_�SCT�cF_UF1__�q
FS�1:�ZCHA�Q�)9�qB(RSD���2x��ޣ�1�0_TW�PR�O����g@EM*0_��V�Tq� �z��DIPҔR�AILAC>��bMFg�LOu��S��9�R`܀��䁟���PR2�%S�a�p!C$�$@=	��FUNC���RIN�`Ԥ�'$fA3RA8 �b ��P#8X0��P#WAR/���#BL�af'�$Az+v}(v(DA`�Q!�(�#z%LD�@��q�#��2Z!ہ�#TI�5�y���$�@RIA��A�2AF��P;A�.3��45�p�r@�MsOI` ��DF_�P�7��Ac�LM��FA��PHRDYJTOR�G͢��fS� �5MU�LSE�P�����J��J������F�AN_ALMLV�V�AWRN	EHA�RDpP�E�Y"2$?SHADOWl���/�?Bc�@w@u�:�_m�ЖAU�`�:�|@O_SBR&�E����JU &�/!�CMPINF��k�D�!�CREGpU��л�i�g� J��Q$;Q$Za4e�O�j���� ��EG0�~���*QAR�����2�q7W� ,�AXE��ROB������d��R�_�]w�SY_��dQU��VS�WWRI8�P=V5 STR����T���EW8�FT�q	kB�`B�P���V,�\����OTO�A8���ARY��3b����B�ƱFI5�ܳ$���Kq1��Sa]�_��S��EU3�zbX�YZ'B�j5�fOFIF��Rbzbnh7`	B��"�d��V�  �cFI� �gq��«�"��_J��6���Fy�$a@dk6��F�qTB)q�2arC� ��DU��DV7�TUR@X
3�uAa�B1X�P��IwFLg�TЀ��7P�p�e�Z�û� W1�8�K��MД�DV����OR!Qy��V#�W3I���2�+�s0�h�à�TNz�OVE����M�  *��C��S��
R��6@ ��*A��W ��<�! � 50�����݀Q�*��������'�S'���E)R��Z!	�E�PD�$�e�A����eH%`t?g�!���!AX�� 6��!Ua���˙ �1˙�`ʚ�`ʚZpʚ@�pʚ��ʚ�ʚ1_� ʖ�0Ǚ�0י�0癮0 ���0��0��0'��0�7��0G�d�X�DEBU-$(!4C����vbAB�����~�9V��, 
#�Y� ?�K�OW�#aW��aW� �aW�ZqW��qW���W���:4fp42���cLA�B�bI�) 6�GR�O� Ir-L��B_ �L��T���`�@ �4�pJ�0�A<�AND����Z���e]�Ay�  ���@~a�ȳ!�ȡ ~`�NT@=!�SERsVE��P� $�p�T Ae�!��PO���K@��-`��p��_�MRAQ� d �� T��e�ERR�r2�00TY2�I��V�`��7�TOQ�����LhP���RJ� � ���D@Q �� p 4��Ԯ�_VA1f����Ԥ��2��!2���D@�p�H��N��$W� �֬q�5VQ��@$���4d0i����OC�!P��  �CO�UNT�Q  ���SHELL_C�FGQ� 5�!pB_BASVCR�SR�AB� �~SSW�!h�1��%�g�2��3��4��5*��6��7��8��[�ROO�0��Y`}`NLQlsAB�úi�ACK4�IN�T�� ��lpa@�0�_cPU�0@�OU�3Ps l��I�����TPFWD_KA1R<ї0�RE�Ę0qPO`�! QUEr�@t��� �r.@_AI@�7�H�{`�D��EzbSEM?Ox0)6��TY*�SO��)�D�I6�s ����b1_sTM��'NRQg�{`E� (�$KEYSWITCH�؎�I��HEupBE�AT�qE:PLE(;��U��F����SNDO_HOM�20O<#REFe�PAR�a���Q�P7�C� O�1�v�O �;rK@0IOCMgt��a��u�lG�HKQ� yDxat�RESUUB���M�"��w�wsFOcRCx�#\�G��OM;P � @��*3~@U�SP9P1��$9P3�4� �0�S�HDD�NP� �B�LOB  �p�SNPX_ASP�w� 0v�ADD��GA$SIZVA�$VA:���0TI�P�'#�A�� � $c�( $�`bRS��"QC7Л&OFRIFHB�S����� NFjODBU�P���%�#�)�ş! �Si�P�� x��SIT�TE��sX��sSGL#1Tab�p&��<3íP$0OSTMT�qU3P&P��VBW��%4SHOyW]5�ASVDTU��� ��A00~Ħ2��7��7���7 �75�96�97*�98�99�9A�9\P �7��7ӱ�6�P�7�CP�3W�pH�91�91�9U1�91�91�91IU1I1 I1-I1:IU1GI1TI1aI1nI2�92�9`@X�9�` @X�9Yp@XI�p@X IU2-I2:I2GI2TI�2aI2nI^�h�93��93�93�93�93��93I3I3 I3�-I3:I3GI3TI3�aI3nI4�94�94��94�94�94�94��94I4I4 I4�-I4:I4GI4TI4�aI4nI5�95�95��95�95�95�95��95I5I5 I5�-I5:I5GI5TI5�aI5nI6�y6�96��96�96�96�96��96I6I6 I6�-I6:I6GI6TI6�aI6nI7�y7�97��97�97�97�97��97I7I7 I7�-I7:I7'�7TI7�aI7nD (�0P.� UPD���"+����
,�0GUN_=C��� `�g�7PUT'�IN\���f<AX|�GO��U
GI��IO_�SCAw�0YSL}OP�� � E% �"#��':'� d�� ʤ�	�P�� �R��F���ID_Lj+�H�I&�I���LE_Xg�V���$d��;SA��� hЂ�?E_BLCK��|M1��D_CPU��@F ��: &�Y�k������b�R ��
�PW"��� 	�L�A�2S�����RJ�FLO5��5���� 8�V��V��t��TBC#�C!��X -$}�LEN`��$}�D�RA��d!$��W_��&�1}�C�2��M�b��4� 3�II� ]���GTOR��}��D��<��� LACEG��p}������ _MA+ p�J� �J�TCVQ�r� �TssڒՈ�� ��� ���JF��$M�ԙ�J���0�)�� ���2/ ~0����ӱ�JK(�V�K:�$B�3,�J�0O�>�JJF�JJN�AAL>�t�F�t��n�4o�5��N1 �ܥ�d�N�y�L��{�� �x�CF/!I�T�v�M?1�"B��NFLIC�# R�EQUIREE�BUOy���$Tx�2�6�z� �x�. ޙ3� \rAPKPR,�C��{�
��{ENs�CLOS� ��S_M� $ ����
�$��A?  o�����  �p���%��������s�VM_�WRK 2 ��� 0  �5��)!L L	#�`������q���_��n�+5UXѠ;M_ ������/�B/T/7I�)$ORk}�5/�/� ?�/-?;?1/r?�?xg/y/�9DYN_�/ �/�/e?O�/6O?O?�]OkOa?�O�O�K��B�SPOSU� 1���� < �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ����
���B~�N�L�MT�����C  �1�IN:�L�0�PRE_EXE]�1��l�.�AT}��J�����LARMRE?COV ��l���DLMDG � "�LM_IOF ��d� *�<�N�`�n������x��ǯح, 
�O����FNGTOL � �K�@A   �4�F���PP��Ng ?�������Handl�ingTool ��� 
V8.2�0P/A2E��x�.p
8815�0���80��33�48966��xi�s
91���p�ra����rod�7DE3���p�c 	F�.0�14i�Y p�FRL�ld3�2���V�X��TIV}�l�J��i�UTO�� ��h�P_CHGAPON=���������L�1	� @��������I��U�7 1  \����>j��4�����VIQ�c߽߇���=�� �{����HG�����HTTHKY�ߚ߬��� ��6�H�Z�l�~��� ���������� �2� D�V�h�z�������
 ������.@R dv����� �*<N`r ���/���/ /&/8/J/\/n/�/�/ �/�/�/�/�/
??"? 4?F?X?j?|?�?�?�? �?�?�?OOO0OBO TOfOxO�O�O�O�O�O �O___,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o �$6HZlu*�TO��uχ�DO_CL�EAN��(��sNM  #��9�K��]�o����_DSP�DRYR�'�HI���@(����%� 7�I�[�m��������ǟ$�MAXZ��t�q�q���X�t����>i�PLUGG���w\�Å�PRC��B�EϋޏП?�OD����(�SEGF��K �������'����p%�7�o���LAP̏ ߮�Ӌ�������ӿ� ��	��-�?�Q�cϨ�TOTAL�0���_USENU̠��� �x���r*�RG_�STRING 1���
�Mڞ�Se�
��_I�TEM1�  n e��0�B�T�f�xߊ� �߮������������,�>�P�b�t�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERRɀ = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat�MH� FaulD�M�AlerW���u���������������� �s���q�h z������� 
.@Rdv�8��.WOR���� �X�//0/B/T/ f/x/�/�/�/�/�/�/��/??,?>?P?b>PO��8�0�q?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�Op�O�O_�2DEV�> ,P�?_S_e_w_�_�_ �_�_�_�_�_oo+o�=oOoaoso�o�o�oPALTD�a��o �o
.@Rdv ��������p�*�<��oGRI� ��t��oN�������ҏ �����,�>�P�b� t���������Ο��b���RD����@�R� d�v���������Я� ����*�<�N�`�r�<���PREG�n�� 0��������,�>� P�b�tφϘϪϼ����������(ߊ��$�ARG_�D ?�	���k���  	�$��	[�]������^�SBN�_CONFIG �kۊ���CI�I_SAVE  �������^�TCE�LLSETUP �j�%  OME�_IO���%M�OV_H!�4�:�R�EP���X�UTOoBACK�
��FRA:\��g �調'`#�9����� ����x�15/1�2/03 07:_34:46�������B�T���x��숄 ����������"�����Pbt��� 5���(: �^p����C �� //$/6/H/'�ׁ  ��_��_\�ATBCKCTL�.TMP DATE.D�l�/�/�/�/.��INI�`���~��MESSAG����!��s�����1OD�E_D&���?E_�O.P0?��PAUS��1!�k� (�7��Κc?�!K*���(��2���� ?���q��)��A��c�/��99���? I�?O  (On�(O:K $OZOHO~OlO�O�Ic4~m0TSK  s=����M�/OUPDT�'0�'dP5XI�S��UNT 1�k��� � 	 �� M|��L<��6 r} ������GP B9� �dy� Y�� �2� ^s �D��b^�_�_GP���n H}� ��R �^ ?��d <���_ ��S�_�_oo@o+o doOoao�o�o�o�o�o �o�o*<'`K �o������ �&��J�5�n�Y��������ȏ���W�)QM[ET�15]Pޏ 7�ڏ[�F��j����� ��ٟğ���!��E����SCRDCFG� 1k�%������@��� ��ȯگ�����"��� E�W�i�{�����
�ÿ .������/�A�S���YԤ�GR.PPQ?�}�j NAN�j�	���z�_ED� 1�t�� 
 �%{-p EDT-k�pb���ߩ1� @�Q-����/����?����.�ߗ�0008�����2H� ������;R<ع�$�k�R}�2�ߢ�2��3��ߩ��߿����7� I�~�1��P��4(�F� ���d��Q�������9���5��d�A�� �������w��6�0T���T ��C���7�� � ��� /gy/����8X/��/$� �/�/3/E/�/i/��!9$?�/q?�/�M?��?�/?�?5?��CR ���<ONO�O�O�?��?qO�?}���NO_�DEL�ϛ�GE_�UNUSE�ϙ�L�AL_OUT ���  gҜ�WD?_ABORT
_{��CPITR_RTN�  /����CPN�ONSTO��nT� ���$CE_�OPTIOkX��ƣPRIA_I�	PnU�P���PFFn�+[ڳ/��Q�_PARAMGPw 1+[�^�g�Qocouo4kC��  �n��`��`���`��`Ș`Ҙ`��`�`�`�  �D�`�`�`��`�d�`�m�a	���bD"p/�`;�pH�`Tpa�`m�pz�`�@ D��p�� D�`/�?���o>ogy��n|�`��`��`�� �C��p��p��p���p��`��`��`���`Ř`ʼpмp֪�pܼp�p�`� �����|;Mv� ���������1�� ŏ׏���I�[�m��� �������-�?�Q������	��i��PHE>�@ONFIGK_���G_PRI 1+[ @���دꯀ��� �2�D�V���K�PAUSPOS s1���S ,]E ������ƿ���Կ�  �
�D�.�T�z�dϞ�ЈϮ���j�O�Q��_%׿QO_MOR�GRP 2l }��0A���r�:� 	 :�R�@� v�dߚ߈�k������� ������2���h�V� ��z��:�L�������
�@�.��c�!݋���?o�o��`���0K���1r�����@�����������PP�½+U�` =Ua�-��k}��:
\�	�0P�N@f��5�Y`�53DB��+Y�I�2)cpmi�dbg[@m:��?(?)�UAp0G�k�`��kP�O�E���`٣����-/�����|�cmg/v/A/�����fe/�/���/?ud1:�/?�7~"DEF ���7)�!c!buf.txt?e?�4 _L64FIXw , � �?�\�?�?�?�?&OO JO\O;O�O�OqO�O�O �O�O�O�O"_4_F_~?�MC�,P � d�_�_�UfS��t]��T�Um����CpBp:�B���kB��XB���B���B���yC=�
;�D�(IC��D�(�VDC�HD?-��Dr<��f�FחF�W�F�NFkNx�F8+/F��Є�	r�4���]��YDǺupT_�;�G����o�oK�# �o�lo~o�Y�oQ< u`�,������;���6g� N=<�	���������أ���ӣ�x��;�C>$<����<��`D��n���Dπ��fE}�π�  Ems��a�πz��C  �F�E��fE���fL��  >�?33 ;��s��n���@s�5ُ@333�.�� A��=L��<#�
�2����/�����~���Q���Q��Ey��� � H����1�9�J;#�H�2�� Z��J�9�Q�e�w��� ������џ���B�� f�=���a�s������� ��ͯ����'�t� s�]��ρ��ϥ���ɿ�ۿ��5�#�v�2R�SMOFST �6>���9T1�PD�E !=�pGX���;�3�U߼O�>TEST024��R7"r��|�| C�pAʀ���U ��!�C�B����b��cC�@i�-�J:d�
-�I_j1�#7�-�T_00PROG %r��%v?��*�T_IN�USER  7e�(�C��KEY_TOBL  ��(����@0	�
�� !�"#$%&'()�*+,-./01�23456789�:;<=>?@A�BC00GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~�������������������������������������������������������������������������������͓���������������������������������耇���������������������t���LCK������STAT`+�_�AUTO_D���%�INDT_ENB� ��П�T2�-�STO�P��SXCh� �2$B� 
 8�
SONY XC�-56L輸�  ��@��ʹt(� АOH�R50K��o�7<��Aff���// �>/P/+/t/ �/a/�/�/�/�/�/�/�?(??L?^?�TR�L��LETE� ��	T_POPU���-�T_QUI�CKMEN�4S�CRE�0B��?kcsc�4�x�0�9��c_�4uUM�0U 1��  <K�% k?gOK�EO�O�O/ÁO �O�O�DF<��_�O_�P_�LStart� SM Comm� %IBSCM�ANS[_�NEn�dxV�@�U�0�_�]U�ser Canc�el�RUCANC�AC� o�L
�RR�eset�BURES oo3_E_�oYo�ko�o�o�o�o�o�@�Zange�GZG_-A�_�ocu L^��������)� ��_��ZVA�G_KONFIG.�RVW)��=�O��؏s�-Datei�eL�%DATEI�1�����E��.� @���d�v�ß�������П"bMacro Step tt�P�MSK_}<��L�Wait Mon�itor3aSHTP�G�L�柫���������ZCYCLE� POW�PPW�D����� DO�W�%	#�_MA�INu�a�%Cb�NUsAL�?�ZCD��#&��C�[�	���������?|(���$DBCO� RI��Ќ5#DBLOV�RD�%�NUML+IM��d����DBPXWORK 1'���ϩ���������DBTB�_1 (7�P��Q���s�DB_A�WAY��GC�P ��=��3�_A!LU��?3��Y�5���$�_DBG 1�)�� ,I��
��#�G�	�ат!��ӆ�$���5�M�� It�B�@��	�OoNTIM�7����)��
)���M?OTNEND����RECORD 1�/�� �D����9��D��D�_��:�lD�0G�O逿��"�����v�����E�XECUTING

 ��	���������D�>EĪ��D:��D��|�Ī� D:k�s��#��.{��w����)�����/��A��u�īg�D)��D��7�ī>!D+N������P��j�ま����Rd���A��h��L��D��D�i���O��DS�d���끾������+/q��w�	�!�D���D��D�����C~hD]������,����B�ONE
 ����"��������h��F#����>/P/ �t/_/��/��B��/ �/�/�/h/?�/?�/ e?w?�?�?
?�?.?�? R?��*/)O;O�?_OJO �?�OOO�O�OtO�O _�O7_�O�Om___�,_�_$_�_H_������_o*o�_No9oGo��oc?�o�o�o;o��TOLERENC@�sBȉ�N�L����CSS_DEVI�CE 10�  üƹWi{ ���������>sLS 11,}�
 E�W�i�{�������Ï��PARAM �2����TuTutR�BT 24,|8���<I�� C��* ���	HR�&��`T�˴���?�g۶�p���  �\  �gI@��˴��A��F�+��p R��Ɏ��f?�B���Ʌ�zɇGă@��\�7�1����q@���Ɇc ��Ɇ���Z�l����� ����Ưد�7�� �|m��C�y�D��C�9��ѰA����A�ffAI���A;33Ad�  A�Ɍ��B�`pѐ��U�̱C>���BffB�;�-��B*갉�ֿ��ҿ�� }<�� �b� K�@ S�D�ɍ)�K�]��� E�sυϗϩϻ���� ��>��'�9�K�]�o� �ߓߥ����������� �#�p�G�Y���3� ���������*��N� 9�r���_ύ������ ������8!3 �Wi����� ��4jAS �w���c�/� 0/B/-/f/Q/�/u/�/ ������/��/�/>? ?'?t?K?]?o?�?�? �?�?�?�?(O�?O#O 5OGOYO�O}O�O�O�O �O�O$_�/H_3_l_W_ �_�_�_�_�_�_�/�O _2o�Oo-o?oQoco �o�o�o�o�o�o�o�o d;M�q� �������N� `��_��o�����̏�� ����&�o/�A�n� E�W���{������ß ՟"����X�/�A�S� ��w���֯������ ���T�+�=������ �����Ͽ��,�� P�b�=�k�}��ρϓ� �Ϸ����������^� 5�Gߔ�k�}ߏߡ߳� �������H��1�C� U�g�y���A�������  ��D�/�h�S����� yϧ�������� R);M_q� ����� %7�[m��� �/}�&//J/5/G/��/k/�/�/�/��$�DCS_CFG �5����!���d�MC:\� L%0?4d.CSV�/��#=��A K3CH
S0z��/#>^?�?.�  ���2�1��?�7� �`i�MU���(RC_�OUT 6�%��!��/�!_F�SI ?I �9#8AOSO eO�O�O�O�O�O�O�O �O__+_=_f_a_s_ �_�_�_�_�_�_�_o o>o9oKo]o�o�o�o �o�o�o�o�o# 5^Yk}��� �����6�1�C� U�~�y�����Ə��ӏ ��	��-�V�Q�c� u������������ �.�)�;�M�v�q��� ������˯ݯ��� %�N�I�[�m������� ��޿ٿ���&�!�3� E�n�i�{ύ϶ϱ��� ��������F�A�S� eߎ߉ߛ߭������� ����+�=�f�a�s� ������������ �>�9�K�]������� ����������# 5^Yk}��� ����61C U~y����� �/	//-/V/Q/c/ u/�/�/�/�/�/�/�/ ?.?)?;?M?v?q?�? �?�?�?�?�?OOO %ONOIO[OmO�O�O�O �O�O�O�O�O&_!_3_ E_n_i_{_�_�_�_�_ �_�_�_ooFoAoSo eo�o�o�o�o�o�o�o �o+=fas �������� �>�9�K�]������� ��Ώɏۏ���#� 5�^�Y�k�}������� ş�����6�1�C� U�~�y�����Ư��ӯ ��	��-�V�Q�c� u������������ �.�)�;�M�v�qσ� �ϾϹ�������� %�N�I�[�mߖߑߣ���$DCS_C_�FSO ?������ P �ߣ���� �"�4�]�X�j�|�� ������������5� 0�B�T�}�x������� ������,U Pbt����� ��-(:Lu p������/  //$/M/H/Z/l/�/ �/�/�/�/�/�/�/%?  ?2?D?m?h?z?�?�? �?�?�?�?�?
OOEO @OROdO�O�O�O�O�O��O�O�O__*_��C/_RPI����@_ �_�_�_X_��|_�_o�0o+o��SGN �7��r`��k��06-JU�L-24 21:�58   ��{`3�-DEZ-15 �07:35�`C`�Ab Ig�aH-ݻa�a5n��`wa���B��?i�ZX�_�o���VERSION �jjV3.�3.2�lEFLO�GIC 18���_  	Gh���Ny��]~0rPROG_ENB  5d�Es�`~sULSE�  cu�u0r_�ACCLIM�v���s��sWR�STJNT�wra���0qMO�|�a�q�/r�INIT �9=z���� �vO�PT_SL ?	�;��
 	Rg575@ch�74m��6n�7n�50��1���#tNy��*wK�TO�  W��o�+vV."�DEX�wdrbC`�)�PATH �AjjA\KJL�TVL41163?0R01\ g�n��-REPASSA�R\�$DHCP�_CLNTID y?vEs Go� ǟ��IAG_G�RP 2>����R�ؑ 	 E�  F,D�E(p �D�5j��B�  =�+�B��C�f�T�CeEC��  C��C�G�SCEZXB��Gm:jf36�2 678901�2345��� � �  A����A�=qA��A�33A��z�A��A���RA���A��ߠ���5j֠Ba@o�  A�`Ap�,�B�A�C�C��`;B45l 5eW��Ba
բ���{�A�ߠ�ߠ�k�����G�Aď\�A��A�Q� 7�� �2�7�F�7�U�U�ߠχ��۠����������A�ffA�۠򠍿�����ÿտ[�_��Z��U�O�
AJ�ߠD۠>�8۠2�,O�&�8�J�\�V�_`��A[��Vk��P۠K
=AE��A?�8��A2��+�
�Ϸ��Ϩ����[��������x�q�j�c��\Q�AT۠L��1�C�U�g�y�[� ��v����Ѧ�-��=�G�I�>8Qy�U�-�8��bq��7�Ŭ}�-�@�;�\���p����m�@*�Ah�а��<��C�<�t�=��P=�hs=��ᗍP-�;��M
��<#�5lÐ��?+ƨC� � <(�U�b �4����A���Y�M�5iA@Ab?5� ���r������:� ������5YkM	?Tz�
�2-��J�G�-�2��C`�-�xC����}�
��/G�{CEY����ɦ4ZH������/��Ҧ�ED � E���D�����m�/  8���Jľ�o�E�s���z�#=�u>�>N�<���?�x=�y����q�*7bD�n3� ���`�o/���/J�/�"5i�E)C�NB�[6�'�/?}/�&??J?5?G?�?D` ����ϧ�?�?�>�?O OD�V��uWO�FO �O�O �rO�O�O�O�O _�O�O_d_v_T_�_ �_6_�_�_�_o�_*o <o�_Ho"o�o�oto�o �oVoHO:% ^I���i����J��>:��6�-� �og�Iw��������� ��	����?�Q��o x��������ҟ���� ���>�)�b�M�_� ���������/�� (�ϯL�7�p�[����� ����ȿ�ٿ���6� !�Zω?�?�?�ϴ��? �����+O=O/�Aߣo e�w��o��]߿��߯� ����+���O�a�?� ���!�k������� �'�����]�o�M�� ��/���g���G��� $J5n�W�� ��	��"Q�C U7�y���Ϗ�� ����-//(f/ Q/�/u/�/�/�/�/�/ �/�/,??P?;?t?_? �?�?�?�?���?O�? O:O%O^OIO�O�O�O qO�O�O�O�O_�O_ H_wωϛϐ_�_���_ �_��/o/ooSo eo��9o�o�o�o�o�o moo�o+=as �o�Y����� �'��K�]�;����� �C/�_ޏɏ��&� �J�y3�X���}��� ������-��1�/ U�g�y������I�ӯ �ǯ	��ŏB���f� Q���u��������Ͽ ��,��<�b�Mφ� qϪ��?�����ϙ�߀�:�%�^�p߂�LU��$DICT_CONFIG ?m���sVzP�egWS����S�TBF_TTS { LT
����VER��xQ�����MAURST�  LT�՜�M_SW_CF��@���ZP��OCoVIEW��A<�����ώ����� ����XR|��#�5�G� Y�k������������ ��x�1CUg y������ �-?Qcu ������/� )/;/M/_/q/�//�/��/�/�/�/?��PM�5�B<�xS��  ����;SCH �2H<�
�yQ�Schedul�e 1 LW ���R䑏9ZP?�?M�HA8�1�?L[=A�4>L�Ͳ2D �?�?�?O"O@OFOXO jO�O�O�O�O�O�O�O �O__0_B_`_f_x_ �_�_�_�_�_�_�_o�TJafeU4ueD5�9m*o �9Dzhg no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x�����@����ҏ�����5=`6�Jeb�t����� ����Ο���	H�V� �)�;�M��?�?���? u�;oMoo����ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ���_o�B�5�G� �7�I�[�m�ߑߣ� ������>����!�3� E�W�i�{������ ��:�����/�A�S� e�w�������S��# 5GYk}��� I����92�?`� r�c��T����ψ ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?��� �?����O(O:OLO ^OpO�O�O�O�O�O�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �&8J\ n�����@ R#�v��?�?�?H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d��?�o ���o�o�o֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tχϘϪϼ� ��������(�:�L� �o���������
�� .�@������ 3. ���6�� ��v�(�:�L�^�p��� ������������  $6HZl~�� ����� 2 D��p�x�ߦ�d߶ ����/"/4/F/ X/k/|/�/�/�/�/�/ �/�/??0?B?T?g? x?�?�?�?�?�?�?�? OO,O��P�O�O�O �O�O�O_ _f��b_ t_�_�����_��_z �V�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��PO8�tO�ODOv� ��������Џ��� �+�<�N�`�r����� ����̟ޟ���'� 8�J�\�n��������� ȯگ쯒O0_b�t��� ������ο�F_�_"�4�F���4��_�_�� �_��:�L�������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ��������^���4� F��V�h�z������� ��������.@ Rdv����� ��*<N` r�����R�� B/T/f/x/�/�/�/�/ �H�??&?�ϒ�c? ��T?�,���?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_>���_/ &/�o(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z���2/�/ ��&�8�J�\�n���@�/(?ԟ�`�5n� @?R?C�v?4��_�_�_ h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτ��_ ����ԏ揤����� ,�>�P�b�t߆ߘ߫� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�򏐟����* <N`��蟢��  �2�V�����ϖ� (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?�� ��x?�������?�?�? �?�?O"O4OFOXOkO |O�O�O�O�O�O�O�O __0_B_T_g_x_�_ �_�_�_�_�_�_oo ,o��p�o�o�o�o�o �o ��bt� �6����� z?�?V?��,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$��?PoX�to�oDo ������̯ޯ��� &�8�K�\�n������� ��ȿڿ����"�4� G�X�j�|ώϠϲ��� ������ߒo0�ߔ� �߸������� �F� B�T�f�������� Z�l�6���������� "�4�F�X�j�|����� ����������0 BTfx���� ��~�0�T�f�$� Vhz����� ��//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?r��BOTO fOxO�O�O�O�O&�h�__&_�z7���� �_��t_,��_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |����>�?� O&O�?6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v�������2O �O"�4�F�X�j�|��� ���O(_����`_r_ Cϖ_4����h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r���Я�� ���į����,�>� P�b�t����������� ����(:L^ p�������  $6HZl� ����//*/</N/�`/ƿϢ/�/�/@Z8 N_ �2�#?V�?���� ��H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ ���_����_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L��p/ԏ��� 
��.�@��/�/���� �� ??�6?ԟ�_�_ v_��,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� �_p�Xϔ���d��Ϩ� ����������&�8� K�\�n߀ߒߤ߶��� �������"�4�G�X� j�|���������� �����P��������� ������ f���BTf�*9�/��ҟ��� �Z�l�6��� 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/?~�0�8?T�f� $�v?�?�?�?�?�?�? �?OO+O<ONO`OrO �O�O�O�O�O�O�O_ _'_8_J_\_n_�_�_ �_�_�_�_�_r�bo to�o�o�o�o�o�o& h"4F���� t:?L??���� ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ^?o��4oFo o6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬ�Ro�o"� 4�F�X�j�|ߎߠ��H����� �10��k\�្� �ϟ��������"� �����j�5�G�Y��� }�������������B 1�Ugy� ���������Ͻ� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�߻�OO 1OCOUOgOyO�O�߻O �O�OYK�_o��R_ ��A_�_e_w_�_�_ �_�_�_*o�_ooro =oOoao�o�o�o�o �o�o�oJ'9� ]��?�?�?�?�?� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E��?�?�Oͯ߯ ���'�9�K��O{������a��$DPM�_SIM 2I����ʱt������C&]Y&Um� � 0�� DϨ�q���RC_CFG Jʵ�!�X� &]���ϸ������ ��5�6ᾰSBL_FAULT K���s�O�GPMSK � &Tb׾�TDI_AG Lʷհ�SQ��UD1�: 678901�2345��xz޻P �����1�C�U�g� y������������X	��Y�۽@��ORECP�ߪ�
�� ~�ܿ�ߴ���������  2DVhz��������9�K�U�MP_OPTIO1N|�[�TR��}�z_�1PMES;�J�UTY_TEM�P  È�33BȱЅ�A�o�UNIT|ׅ��Y�N_BRK Mlʹg�EDðZE|��'t�c�x�TA�T��EMGDI��[��NC#1Nʻ ��X/K/&^u�&[d���/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>COUOgOyO �I�!�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo �J<OFoXojo|o�O�o �o�o�o�o�o0 BTfx���� �����4o>�P� b�t��o������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �,��H�Z�l���|� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
�$�6�@� R�d�ϐ��ϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��.�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������&�0 BTf����� ���,>P bt������ �/(/:/L/^/x j/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?/O 2ODOVOp/�/�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_O O*o<oNo`o zO�o�o�o�o�o�o�o &8J\n� ������foo "�4�F�X�ro|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� j�t���������ί� ���(�:�L�^�p� ��������ʿܿ�� ��$�6�H�b�X�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ������ ���.�@� ��l�v������� ������*�<�N�`� r��������������� 
�&8Jd�n� ������� "4FXj|�� ����//0/ B/\f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �OO(O:OT/FOpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�?�_o o 2oLO^Ohozo�o�o�o �o�o�o�o
.@ Rdv����� �_�_��*�<�Vo`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟB����� "�4�N�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�F�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������ � �$�>�4�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
��H� Rdv����� ��*<N` r��������� //&/@J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?��?�?OO8/ BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�?�_ �_oo0O"oLo^opo �o�o�o�o�o�o�o  $6HZl~� ���_����(o :oD�V�h�z������� ԏ���
��.�@� R�d�v��������� �����2�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� �����Пڿ���� *�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮�ȿ �������"�,�>�P� b�t��������� ����(�:�L�^�p� �������߮�����  �6HZl~� ������  2DVhz����� �$ENETM�ODE 1O��  
����������RROR_PRO/G %�%��:/�G)%TABLE  �%�/�/�/��'"SEV_NU�M �  ���� !_AU�TO_ENB  q%�$_NO�!� P���"�  *�20�20�20�20� +10K?]?o?4HIS�#����;_ALM 1Q.� ���2<��+p?�?�?O"O4O�FOt?_OUT_P�UT 2R�= G @ٌ7���$_�".0  �01���J�TCP_VE/R !�!2/VO�$EXTLOG_7REQ�6�9S�SIZ_TSTK�;Y 5�RTOoL  ��Dz�2��A T_BW�D�@xP�&�Q-W_D�I�Q S�4�����VSTE�P�_�_��POP_�DO]_�FACTORY_TUN�7�d%iDR_GRP� 1T�  �d 	�O|o�m`��[���N�8�T&�hB�( ����fmc�o�mm`�B��xCD'��C'��B��)�B���C���mA�pB8L�0B+	A���}A�dEA�����n$y��o�o��n�Q��TA�^4m����??�A;����0|�8V}B��A�� gA��A���A���m����R�Ҹ�����y�������A�������m?�x�AW��A5D�?����?���?6���Kz
 Gm��Zq�qhqAÌU�K�2�aL E��  F,DG�E�(pO�DE�4�D � E��o�D��xw�m��mC��N���B�ƈ���m@UUU��U��o�=�?�� E�@�����mOHcGP{8�L�uS@�K�y
�~"�\����:G:���9{������m� @ �[h'����9��.4����|ԏ�o�o00%U6�j	��o0�ۏT� ?�x�c�������ү�� �����>�O��pO� u�$���9�����ڿſ ���"���X�C�|� gϠϋ��ϯ������� �͟?������%� ���߫��������,� �P�b�M��q��Y� ��}������:�%� ^�I�[���������� �� ��$6!ZE ~-ߟQ�c�u�s� o D/hS� ������
/�� ./@/���v/a/�/�/ �/�/�/�/�/??<? '?`?r?]?�?�?�?�?��?\JFEATUROE U�U�P	a�Handl�ingTool �'E ally�English �Dictiona�ry-A, Pa�Multi L�anguage �(GRMN) t�\ir4D �St@ard'F � prodA�nalog I/�OzG  VLOA��Agle Shi{ftzHl.pc�@�uto Soft�ware Upd�ate  \pk�4�Cmatic �Backup+Ci�rpk�Agr�ound Edi�t @-A�@uC_amera�@F�I��@DPnrRnd�Im�C)E�@Po�mmon cal_ib UI S �@Έ@ConQSPMonitor,B�@�@�kPtr%@Reli�ab�@,Bduct�Data A�cquisoS,BA�D p�Piagn�os�A�A*D
PC�V�Pocument Viewe{R�.@wc.�Qual� Check S_afety[Q �P�l@Enhanceod Us�PFrP�.@ENDI5@xt�. DIO kPf�i�T *`F-ben]d`ErrzPL�R�dTKfgs  ck�ToIcr�@3` B�WD*DINT �FCTN Menu`v�S�AM@�`�TP In�`fa�c�e{`t\j�G Pp Mask� Exc`_@�EH�T�`Proxy �Sv�T�A�QHig�h-Spe`Ski;TdPcs@�P7`�mmunic�@o�ns.@�P\)qur��`�`�I.P�`�A�bc�onnect 2�EWIncr�`st�r�P�Vcsge�KAREL C�md.XG�e�sRu�n-Ti$`Envz�WK�`el +�@]s�@S/W-A�P�Licens9e�S�Vetw�PZ`�Book(Sys�tem)*D  � Q@ACROs,~r/Offse�@�HTMH7`�@J��@n�gQ@echSto�p�atpp�RPsi�Q@iUb�K p.f�@Mix`�@�@'G�t`Q@od�@wi�tchzH93 R豁pR�Q.E� R8{08͆OptmڈrPJ͆�`fil�VGt I,`τ�@gOw� 0\t�PSB-T��`
SIPCM fsun�w�cF OY��v�pRRegi�r�=p�qGaPri�PF>`� ELSE���@Num Sell�  oadx���"` Adju-p*DN@�l@˕�J \j76�tatu��Xx˕��Y  F`�`RDM� Robot>@s�coveGA imN�Remj�7anqG� !b?�Serv�o7`��,B!��?SNPX b�rzH�596�`�CLib9rFC۔H55��@A {���〙`��o�p�t�`ssagI� ~�aTCP �C�8�}K��/I�m 1|�p��MILIB!��.vrLP�`Firm�B'Gj7á�`�b'AccP	U
��Q��TXJ��55�T�eln8�"�55 a(��$A4�h�I)�`�Torqu�@im�ulayQQ tp�h�@Tou��Pa��q'GP�� P�Qփ&��`ev.  i��USB por[t SPiPN`a�P� P
!1�neOxcep��Y�n�S� 9 R�i'G ["L�`VCWQr8r/rp�ڰ"���P��\�����@�ı��T��SP� CSUI��hcl�P��XC��MA,`?Web Pl�.�ER�`�y�O{�p̀�/��`d�Qz`R��?�<ZC�@e�Gri}dD�play BA`e���D�QJ�iR���.qJ���ԍ�AAV�M��IO`pNa�PAxy`,B77����-A�TXPL�+CHC�SB9�-2000�iB/210 V �b\��Ascii�aΒLŐ�P��L�c�UplŐ'G���A��f�`opPBA 0����A�qW�����1�`C�E�`rkJ�g R=7PPRUT�����LQRT/KeybowAMan^@v�:���PC�Pl sd�b�y E-c�Uol�:@qQGuwF|�C�P��@�@b�QkPss@tzN@t�� td\$�Eo�prE�s@�f ���LQyc�@�r��or�i`��P�PCS Jo��sc`����@0��a�Blu 4e��P�H��<ZF�,`D�@i�n N#ay�.�5�LPDy���if=i�S 10i�`f�DG@�p/�cUb�Outpu�B0�ࠃ`����imiz��tym��KfAxis7a��Q �����fm��s޹�  MS��FR-L�am� ��P@HMI Dev�p (��� ␠P�a�ΐ��PM�h77�2�p.qnn/Cr֐oޑ�@J��x�o� #1��u��773.=��dЃZqKRD��O���Qb�d��C�o�qTXY�ROFINET�J "AM0�d��Dp�GRAM/J�OG OJ����@ �! d�Passw�ol�i�R�`5!th�����8�SN�`C�li�Q#XM ��SP�EED OUTP`���c`�� RHiĺ�s=e801DpVAGn�r��2"�!`vogi 7��BL$�#z��3^.WeavI��~*��V��64MB D <Z� Ġk2wFROs;802DpwArcҐviszS��*Auxx�J&Ce�ll�L6�9��OTsIh�1(FM�@�<c݅h]s�5�@p�  m��7ty�@��@r2�@����(9���� �� p1`۔I���w�.�/s��PR�� 20P��Q7� e�@`�LR�ZvE% �Pu+�DDf?�x��Pq`@5L fT1G�T8���w40� ���D�s���,���t�BOP!T��pQ�SN`�`�cu�[Re� �p��Syn.(RS�S)$QlU�quiry`		 0��?������ @8�t�
�Qe�stSm0t-ES1S�) ՠteHPWy�S7@��miLjECS�p�a_�N�h681؉$r'�dib� LJ���P cR��q��<p�| iA/l��a71{ap��=��!{a�Z� END  ��d�pn���fd ->�#V8.x I��(��!EMZ$�EQ� ñ����LF�REU �e��d@a1 �#�s\0� �+ �� 8�whe?n arg j�!����͡CD�tiBp*=�Qk�͡u8s}d R.Skif��WF,� BCK �TsAb�v!a�un9g�pϠo�!r�j�P�!1�q68���I�Q�A F�`b.�Tig/Td�(C�� ix up�� }l�bof GOس�To f��G�p�Q�m�psfmn$�p�s�tQ� �:��-PS-s�r�pL|�@�Aff.a.d �S.PN:FW-CHK JG"��� ��\cdc�CD:��SSTE=P̢BWD <􏀿.Er.af� �8xVag_C.2l�j ��tseJ�� �Iss8` iq��+P.Alloc.Mem.쀛k�329P��� I�����w .K[�l Va�r.Scr &�O�����FB_C�MB�lar��MNqSࠏ�I�wr.�!�FUNC-Mx�R9`���	s � S��˓k�n.sMP 6���Z�cmd.e�r.-Pdl.�Pr�p��aEC#rign�Ǳ�& f� }�TSHELL He�beat���Noށ.On/��w.SRVO ?!���t,�9�m�� aw���6��GunM.D�O.@!.Gen.�A R71l���?��.scrn fr�eeze q�P381+Invn9`ig.��ch�p�eldpŁx ABC&"g�p~�X '!�.d��.uP�p.���ar gex.�4�.��.ab�d PGPX  �R`�k�.��spd�dѐ4����p�� �P}й�۳3wp0�տ��F�r��Rd��/�E�C)��sg�.E�;�!aσ� �Anl}ϟ�R788�ϻä0W�����<����anlg���"�`\	�+ӲPp%�GӁIS�A�c�Ur^��
xY�yߛ�8 J6����(Lin��S��<����o\aw��ϐ��ӿC��Pk=��e�coY�{�wmle�u��MH Dϳ�4g8 H���MH�����Tِ���d "yF�#�\mht�p3�b�:�[�"AP�w�htot���B��ί�ETU����ol�$�.������l �E=�5o�c�sQ�)�;���
�4�545`�:�I�p�����H57�4��J�2���fAa����`��j� ��cenl��̨���H50��INT/��`-/�ķ�I/`k#a�f/�z�55���-��/�#9��/'52�/�0K��J?g"MN�/�50� �4�r~?�2Z�!�?��u�4J6_P�?�2���?t42�+D&0M`%O;ūpBO� "@O0��azO�Bic���O�#0�/81�O�CpJ�O_']��"_�Ӷ�f8�ENY_lo� rϼ?-�_�1�O��AR/��*�o#bx�P�o��! ���- 	VUo��Roo8�ϯdg2 J�o��Vi����A0�o�Ds_�.�f ��ib���CLo/�_2�O��Mp��;?�}vm\#cv��Yt�T�sT��Egnai�`�?]�����O�taX_`N_4/a���a.@���cb_-����Ő�e�;�a�a���bsi��w��ޡ ���dӟ1Vig|?�l/~/��r+�=���a�S�𯗟y
n'�9�F��H�|�G�nP��gί��ѿ  ѐͿ�� A��531l~wO��O R=ϫ�RS�?�� F�6E09  ��W�o�_P��dmTo¿H�Z�X/u߁ ��U�0����A����/��_�SEN9D���3 RX�r6���efJ9�Ϣ�AC�4��P�_��mnm��~��.�x���CR�L�*�\sf�v61���j�/�6Y@i���	fK�	�j<��ߌ����ND���1p�f���fe(F�?k�3)�e�DB/t�f���ZO�W "H�Og10F��fe"L��5, �o�t\h a���}���3T3tr��^�h6h�J�p.z��ʕ
I%/����n�hm��buD1E��?��F ���V96��4G.$`j_��rl���/��0u?p;��/�?YSC (?:?#Ff��_�e��d9O+�H?�u74TO�D7 ( ?�����	��O^�L  feI	n\/�gJ5_�onOΏVJ51�O*VI)�_�Dsfm�_/E�_b��e8�~_xO48�O&"ad$��I@/&��mn�o�c� 4Z!3 j�o#sioF_&X_59�?3t8.o ingI7�^p�o��t��|��5P���! Lo�w(B�8O����PxE��σ���}� �o�Oȗ����l_��/"/��a� nitL�/�Epl4_��!
��on|�Ƈ��e3 G�JETX�:9K���674=����N #`�n�gcr���/ߥ~u�ɯ{d.p̔���da���74 �ﾯ`�r�HG�q��2.p�vu����/���\���  u:�2��c.p��21k��3"�ݱOR78"�= P��0�J614���(�ATUP  :�OY�545��Y��6��s'�VCAM�/�CRI��=�CU3IF��Y�28O���wNRE� t.vA�p��_ �`A�SCHO@~��DOCVO�{ -��DCSU� p��J60^��0��oEIOCw�NT��S54"�i�2��9��� Ski�SET�w�q���1�J7��9�21@�MASK � K207P�RXY�s��7�9��OCO{p�@1�3��ҵáQ{pkmaY�Q�m�39�s����kcklLC�HN�=�OPL�G�A�J50~�r@I�HCR�PE�IЃCSj��`l��Ђ�K�AR��J55^�rwt FI�DSWo3@�q����q�f`nI�PRr����f����R��aU�CM���ӡP ^�j�T���f�9�1�v���L1�f�����v�2;09��PRS*�́rY�9J�V�FRD��<��|�RMCN����93R�n�|�SNB�A�@1\k��HL]B��ME"��M���������q�2R�in�'�TCj�1�TMI!LC���A®�p= )�cPAб�A�TX�P7krc)�EL��Y���Ү�Y!Y�8E�rc�fX�C�.��Y�95����95f�f.v�|�UECN���UFqR����X�VCC���v \�VCO��1.�fL�VIP.�73�5.��SUIpL� U��XФ��WEBj��1�T���	���2��g J�T�CG��s�IG��I]% PGS�3% RC.�I�s���\at��H89v�8�U1�X��@��H60.�Q�l�R7��]�Rx��t�69����9����� �"Cp�61���J8��0Fp��v��q��7R�j670�3^^�"FSGY�8^���1��6~���HA�4Ĳ�΀X�~�m�55�v�ftp$ J56�������R5��7�%��R7��tun&0�98v���5e�UĻ82��sgt<�5����/����0.�7�0\$ R55~�9�79��J76R�O��0���573��J�96ѱ���"��g���.�T"0�6YFD> ��4.�)p� J�ℊ�p�9����� ��57 �5�A��~�D���\� ��^�b�� ]�����в�I�����V�5��tdf�����^���9ѵ�D;06^�mch��"pm�� ����SVMr�7men��LIr��8�v��CMSF�V"�� j���TY��6�I�CTOj�U���.�sgm��5�����NN��K0f�mkuN8�ORS���%8R��$8��lwEX�T6 ��F��I#OP�I6 t� ����/�R�6!!� ��PRQ I ��8L���Sd2�w�2f�I�ETS�6 U�SLM*�sveg�!6i��52^�x�� ��iase)��OA� �)�RA4N�&�3��VA����IPN6H@.�=�E�ZE�0�  UPD�~�%�U�MC~�1�P1I�3E0}�3�@ "��@~���@^����@�&�@����X�P1"�
��B.�9� �Bf��T2"�I#�@���al'��@����P2Q �B��n�`�7P�.��6R~�tol���P2}��P22v�#P2��m�sP&7P~�kse��sP�?�P24^�Fpl�7P`^���P����S3U�wkks��P27v� � ���P���B��óP3���P4�1h�k��P5}�P5�iQP5I�a�P3y3��gkdf=e��������3J���U��sgkt=e2 D=e�����
=eI����k=e1"������ ��������>��f5B ��ABVe��e��e>� ��qB�e~A��1����2 ���2����e��e� ���>eV!�e�A���B ���ҶeJ!��tQ�f � �e2Q��=R�uJQ��hst.Ev�v `��m��e�!��ft�P �v�g�R�����������n����4$�� � =e"Z�<fak�9�v5�o orcm=e"CC�U�܇cc�f���d9��f�� ���¶e]��g/`�:hm���hlo����9�k 
�T�֟�}y����!H0	�yfk�weyoY���ve����}���unp<f�z���fsub�z�c�fccce�@+��fE�W�i�{�v��������Ğv����뛌�iY�
!s����� �Di�����f Rn�vT "(�58��v� �vcs/ "�: ag˗9251"����f26' �fr���E^j�4ᨖ� "DG�/�ad1g8v��on ��,vM�߄vr��q�?d3se��:�di���r��!�e�d -=eAe	�yf���fN-��f82 vs�I�[�m�8v�Ϸel�Ϯ��ǋsl8vG��T���S	T��/�l�0�B��0f�L���p�dtHf����dg��b�����'�8������dju8v{�41�g�w��4�f5�1�v2����n��r�o�fstK�natz�f0��  �=e������PG�`onSpox�, �Pȫn�OFTt|�bp�feqi�f���alu�f"W�E��͌8vsweq���E�7`tpȦu� "p�&V�n�w�vK"�v��on�f�vz��ui��A�PF@�΀�s��f�tp�f����TP������bw8vI��H���&f��-\��3OT#/5-dvG/Y/�k'K93P�/�kq9P�/�/ "K����/�  H55
P�!I1!IK946!I�!I=�a!I�1!I�Q!I�3@!IA!I9!!I�05!I q�!Ii!�J�0!I9a!I��0PJ�!IaqJ"SAC!IY11J�!IP�  !Iua�J�!I�qZ��!I���Z�!Iin.@J�_we�_�_%V�� 1_X�p�_�Yu�J]_o[=o?[ld_o�[_Kpo�_�_#Ghomj<)�!Ig\ff!IU��1O#G��O#Gaxtd�O�O�o�oa��o�Y�ax�o'��4ASyswas��n�#��ztp�Jt}1Q�h��FGMQO�cG� �J-^h5 ZA�R"�k�0!Inrg�j-M510�O_ės " �-�0\s`zpyaJ��JMNI��Hfmn��)1Z]����NJP"q�cGm#nm�Z�M^�0�~_�[t ���1���qOÏEWT0Z�m�����椧PD �]MpsyȠ���dFFί�Zrl`��0��0�FRA� �`zm��* E����cer�ZM�_�RSo�1�y������Ɵc� `��?K��CLPZ��}tpsZ]�o�P3MA���Ims�J����n���ym���#π5�7�Y�낀�}��G�RD��]B��bd !�-R"�]�"�DN0!��"�odt`�-B"�@-�"�=�r�P"�r^� "�-�"���"���"�����S��"��r"�n�i�1�C��EM_�!�emd������������� �
ss�p
t I)q"�awsde!� !  �� us@
rsal�!�!
IAR8=31din$�<m� Par��bޢ\srg�F { !�
! s��Serv�IF �O�37 R�Lwoad�rvo��I)o�R�de�f.�s+! mi*G C���0*�8- !+�Тng =M�E, P����A�gco��pLN�migp*~F�*�� ��q�=0�f.�s*-��0e�NmDO;fd�+ -�+�ive��²)69�1!:RIN�701�pti*���2I} �+j`:j703�* OpJ�?Oz!K3�set,!?��O�?��+M� �:d�np*ER J�1� R6ZT_+ (�MI�voi@* �"�+��?$H6�*g{.f@*Jog��R52��che�@*^  j�r�_Wogހ*link�k sI/Q_#H J5A;�P0* J8�j/O�,���B)cl�*v�
�J~`�*ppr�x�Jro0z�o�k J68o��B(�P :]�r/�(mPj��oSimp�te�+/R609�[L�z�,�o�ZtoPjspa*�tch�Jth *A�ST kHST�*7[94�zin�T���a?Sta *����Aϋ���b��_��5p.pJCP�|5y8�J�ModbAO�SObt�;��+P�RO [ �O"�93q0�;�/:30\0�_�+FSW�}�o�h9pZam����*�t\j�p J�? ư�Co/�]]=-olp/�N���=8\gpJ��0���RCo��e��Np�}_i0*VM`���_�[�0 j92o��P�ceN�:�M~Pv0:(N?+ WC�On�)dnw�EN�:���- L�I/�F kJ5��r w�:ar��rj�?�}@�cm�n# a0�M=.�0�����U�g�)�c�p* j6�TorP_R�D)�=oOkM�CR HfA� H�j�=1\�;�=�@�*^�@*h f�z-@��82 (a*r :������p�����P:982�*�0�0�B��'0_�S@q�����������0���P:580�*1�\ ;pa��j����5����We�mOk�m�4�\n�-A���8c04 j΀ �usO��-�\�ڍ�a*n �p:�M���ZJ9ϫi M !
mq�M`q�p�z-j~,moo� �����@��i7�J�� zm��/cυ( l6�
H�5;806 �M�5�4_�nN�`�cz\�P���  �STD��LACNGK0-�1Em�C%E<��%E671%Em��%E (SemFChEa%Et��%E�� %EAj]@%EM�%E��6IG!�F- wO)A-%E�Cmp%EJ�HM�%Egw SV%Eo H�F�>�PIGPHF�!%Eh��p�H�F���Fn�mFf3unIO�83`OrC=t%Ectio�F=0x%Em�%E83\s%E�q�G83�H8�FD{ j%EutpumF,] �G19UF9/@"U=�%E(`!V%`mF��x%E�@pf846\%E�m�mFj84%Gg wM90%EHiOpg�2hm!%E�%E00iA%Ept,�F�%E<͑%Em94l%E���f>��fZ_l_~XIn9t�FQI758�_
�FXfrfaPV�_'Cg58\Tv�k75�o��FL-�O;�-��o��k-ne�V=1�RBT
r�P_�9�\f0p_��S_��p9�OPTN�B5ލ�Safe��by� F��QB��586<@��6q��=љ��� �э�]��������!���r4��]r��irx��}R�� Tri������25 H��P�RA����o�Q��rD6Q~�C��NQ��gRq@��]!���q����O���!A�� ��F�Q��j{62��! ma��w- P��napȆF��96�iBZ�(;�p���/�%�DPN)@� �е�I���U���PClu�����B��7҂��݃ۤa��1����������pΒ���Ҭ�P�IZ�]�������N��R754�k�I�0�bskl�����]��萷�1^���sr�t	s/A��D]�妕����J91���!ƺ�C�USa���g�itp�l�g��g���g�sd9m�g�Sys<@gü���R SMe�J737��Qf�P��#DsK�g���Ie���Ne�\sy(���s���menueŎ����Dat0�g�etw8��Ň�740��i�ng� (DT�.bO���Pare�9rf�Er���Βg�=�g�I�s�n�s� Upe�m�g�s07{���R72m�y9ǁg�4 R8���7�pR"m�E�7 �(AE�j�,E�>0
tE�f�dE�in\P�<�RRascbE��B�R- TOE�rt�s�%�R�RD�R61�7E�01��j�R6���609��1�j�TQS]�fo`R�BR��B6�qs4���U�!� cnE�Cont�E�prE�m�R56� JE啲RJ75M6E�lNO�Rc5P�E�q��"q��nsv�E�E� 5�� E�bdmr th��iv��ْ��55���0�����58��J���88,��"OB��bO穒`�淐^�NQB$mb�����v�B$h848rE�2�a�� 48s�lUbB&��9 E��H612E�w� (��250F]Y�j�Lf�
\s���N���i�h61��2090��R H����uL�3��B/1ybB$�b�\]�b��ae�GK� I/��E	79�P�$iBj�(EG]e��/$*�gd\gY�#�gd��cy� C�'T9r�p 22�煒��4���4yclX&a#ck8�/?5t8&��$����U��er�|����4�H��CV�T��KL�� PH`(���L���`90�c30�8>�^94ǀ�^M����:E3 ��  ]$C�L\����9���$]Zq@]9M�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r�������຿̿޿��99�G����$FE�AT_DEMO �U�@�A�;�   �N�D� Vσ�zόϹϰ����� ������I�@�R�� v߈ߵ߬߾������� ��E�<�N�{�r�� ����������
�� A�8�J�w�n������� ��������=4 Fsj|���� ��90Bo fx������ �/5/,/>/k/b/t/ �/�/�/�/�/�/�/? 1?(?:?g?^?p?�?�? �?�?�?�?�? O-O$O 6OcOZOlO�O�O�O�O �O�O�O�O)_ _2___ V_h_�_�_�_�_�_�_ �_�_%oo.o[oRodo �o�o�o�o�o�o�o�o !*WN`�� �������� &�S�J�\��������� ��ȏ����"�O� F�X���|�������ğ ޟ����K�B�T� ��x���������گ� ���G�>�P�}�t� ��������ֿ��� �C�:�L�y�pςϯ� �ϸ�����	� ��?� 6�H�u�l�~߫ߢߴ� ��������;�2�D� q�h�z�������� ���
�7�.�@�m�d� v��������������� 3*<i`r� ������/ &8e\n��� �����+/"/4/ a/X/j/�/�/�/�/�/ �/�/�/'??0?]?T? f?�?�?�?�?�?�?�? �?#OO,OYOPObO�O �O�O�O�O�O�O�O_ _(_U_L_^_�_�_�_ �_�_�_�_�_oo$o QoHoZo�o~o�o�o�o �o�o�o MD V�z����� ��
��I�@�R�� v�������ُЏ�� ��E�<�N�{�r��� ����՟̟ޟ��� A�8�J�w�n������� ѯȯگ����=�4� F�s�j�|�����ͿĿ ֿ����9�0�B�o� f�xϒϜ��������� ���5�,�>�k�b�t� �ߘ��߼�������� 1�(�:�g�^�p��� ��������� �-�$� 6�c�Z�l��������� ��������) 2_ Vh������ ��%.[Rd ~������� !//*/W/N/`/z/�/ �/�/�/�/�/�/?? &?S?J?\?v?�?�?�? �?�?�?�?OO"OOO FOXOrO|O�O�O�O�O �O�O___K_B_T_ n_x_�_�_�_�_�_�_ oooGo>oPojoto �o�o�o�o�o�o C:Lfp�� ����	� ��?� 6�H�b�l�������Ϗ Ə؏����;�2�D� ^�h�������˟ԟ ���
�7�.�@�Z�d� ������ǯ��Я���� �3�*�<�V�`����� ��ÿ��̿����/� &�8�R�\ωπϒϿ� ����������+�"�4� N�X߅�|ߎ߻߲��� ������'��0�J�T� ��x���������� ��#��,�F�P�}�t� �������������� (BLyp�� �����$ >Hul~��� ���// /:/D/ q/h/z/�/�/�/�/�/ �/?
??6?@?m?d? v?�?�?�?�?�?�?O|O2M  )H HOZOlO~O�O�O�O�O �O�O�O_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o *<N`r�� �������&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���� (�:�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ������0�  1�,�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\�n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿��(�&�7�:�-�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZl~� ������� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�?�OO&O8I�$FE�AT_DEMOIoN  :D�h@��3@PDINDE�X]KlA�P@IL�ECOMP V�����A�kBKE�@SETUPo2 W�E�B?�  N �A�C�_AP2BCK �1X�I  ��)MAKRO900.TP:G_3@#%�E_?Z&_c_D:G�E1__UT1]_C_�_�_y\2�_�_UTA2�_�_1onoy\3ooUT3eoKo�o�oyU@9H�lJ3@�@ 8u�(��^ ���)��M��q� �����6�ˏZ�ď� ��%���6�[���� ����D�ٟh������ 3�W��P������ @�¯�v����/�A� Яe�������*���N� �r�ܿϨ�=�̿N� s�ϗ�&ϻ���\��� ���'߶�K���o��� hߥ�4���X����ߎ� #��G�Y���}��� ��B���f������1�t�K�@P�O 2�@*.VR:���RP*����#S����yU�n�PC��RQFR6:��4��X��T|@|�y�_@xI�xV*.Fq�D%Q	�<�<`�STM ��Д" ��RPi�Pendant �Panel��H �/�/�Pi/�
GIFs/�/��/F/8X/�/�
JPG�/!?��?�/�/q?��JS�{?�?RP73�?O?%�
JavaScrgipt�?�/CS�?�(O�O�? %C�ascading� Style S�heetsTO~P
�ARGNAME.SDT�O�l�\�O�UO�1�D�O�O	PA�NEL1�O2_%@�_[_��_2P_��_EW�_a_s_oZ3 �_:oEW(o�_�_�oZ4Xo�oEW�oio{o~�DSHELLp�A %+rCm�����GZG_MENUE0-O�u�q����EEINGAB�J�%3�K�L������vSUMM_�VAG.D>?�O:ķ�������yTP?E_STAT:���;�S�y�����E;�INS.XM[ҏ�@����o�aCusto�m Toolba�r ��yPASSW�ORD�oU�FR�S:\C�� %�Password Config����G�CONF1 ��]��Aǯ����,��y�EXTSERVO C�U�K�c�������U?IO_SET|��%�AϿ	���4ϣy�VWEMZROU S�e�S�kϑ��ϼ�K�AGV�UP[�m��� �ϙ��@���d�߈� �����M����߃�� ��<�N���r���%� ����[�����&��� J���n������3��� ��i�����"��/X ��|��A�e ��0�Tf� ��=��s/ �,/>/�b/��/�/ '/�/K/�/�/�/?�/ :?�/G?p?�/�?#?�? �?Y?�?}?O$O�?HO �?lO~OO�O1O�OUO �O�O�O _�OD_V_�O z_	_�_�_?_�_c_�_ 
o�_.o�_Ro�__o�o o�o;o�o�oqo�o *<�o`�o��% �I�m���8� �\�n����!���ȏ�W��{��"��$F�ILE_D�� 1�X������ ( ��)
SUMMAR�Y.DG#��MD�:W���s�Di�ag Summa�ry����
��SLOG��p���۟������sole l�o����TPACC�N�v�%^������TP Accou�ntin=���F�R6:IPKDMOP.ZI
�j�
�� �����Excep�tion$�ի��MEMCHECK���������/�Mem�ory Data����� �)>��HADOW�������)ϸ�Shad�ow Chang�es,�ߴ�O�)	FTP���χ����1�mment� TBD��ܷ\+��)ETHERNET��͎f���3����Ethern�et 3�figu�raC�����DCSVRF�ϊϜϵ߸��%z� verify all���cĐe�u�DIF�F�ߓߥ�:ﹰ%=��diff<���|f�z�CHGD11�8�*�� Q�����9�}�2����C� ��j���G�D39� �2��� �Y���}�UPDATES. ��Ћ?FRS:\L�7�Update?s ListL͛�PSRBWLD.CM{ό7�N�0�PS_ROBO�WEL��g�:SM�p�)��M��/_Email��aïcį���Տ� ��� /��$/�H/Z/ �~//�/�/C/�/g/ �/?�/2?�/V?�/c? �??�???�?�?u?
O �?.O@O�?dO�?�O�O )O�OMO�OqO�O_�O <_�O`_r__�_%_�_ �_[_�__o&o�_Jo �_no�_{o�o3o�oWo �o�o�o"�oFX�o |��A�e� ��0��T��x��� ���=�ҏ�s���� ,�>�͏b�񏆟��� ��K���o�����:� ɟ^�p�����#���ʯ Y��}�����H�ׯ l�������1�ƿU�� ���� ϯ�D�V��z� 	Ϟ�-ϫ���c��χ� �.߽�R���v߈����;������$FI�LE_7 PRF �����������MDON�LY 1X�� 
 �q�H�� l��y��k���U��� ��� ���D�V���z� 	�����?���c����� .��R��v� �;��q�* <�`���� I�m//�8/� \/n/��/!/�/�/W/��/{/?�/?F?��VISBCK#��2�*.VDM?�?0�FR:\f0ION\DATA\�?�)20Visi�on VD file�?�/OO3?AO +?eO�?vO�O*O�ONO �O�O�O_�O=_�O�O s__�_�_d_�_\_�_ �_o'o�_Ko�_oo�o o�o4o�oXojo�o�o #5�oY�o}� �B�f���1���U�������MR�2_GRP 1Y���C4  ;B�r�	 .�ҏ��πE�� E��@�������πOH�cGP&�L��uS.�K�y
��?�J���π:G{:�r�9{��~���A�  ����B�H̃C��NƕB'�ƈҕ��΄����π@UUU�U�U��S�΁>t��>S��=��h=���>�߂=��;b��B�:{eg:�s�X:+N:I9��2���V�����̃E�  F�,D�E(p�D�����0E��5�D��=��<Əd���� ���������οϊ� ��:���_���nπ� �Ϥ��������%�� 5�[�F��jߣߎ��� J�\��߀�!��E�0� U�{�f��"���F��� ������A�,�e�P� u������������� ��+(a�߂� d�����' ��������� �����#//G/ 2/k/V/h/�/�/�/�/��/��_CFG =Z��T �/5?�G?Y?��NO ����F17�3�0h?RM_CHKTYP  0��r���00��1O=M�0_MIN�0r�W���0��X���SSB3[��_ �
D�e; C)O8K��TP�_DEF_OW � m���PGIR�COM�0aO��UN�C_SETUP  ��%O�O�O�O���GENOVRD_DO�6}�mEU�THR�6 dUd�T_ENB�O ^PRAVC��\�7�0 ���_�/��_�_|O�_� �_(o�_Lo^o�_mo oo�oyo�o�o�o�o $�oHZ�o~�h�3ydQO�@1b���r��eB�8��^���
��';�.�N���F��F�3G�R�'	���ß	�Ær��DFr�t >p0��x����B�80P��B���r�	�y���!�&���"�D�F�x��������k� ɏ珑����1\�>� �:�\�^�����˯Ɵ@����ܯ ��At� V�'�R�t�v���ѿ��ޯ����OGRSMTkScrY�p�0w��m�x��$HOST�C21d�y�0�IQa}U@k���A��k1�72.26.29o.230��e�� *�<�N�`�n�e�ϒ��߶������� e	�cfg_fanuc���.�@�R�b�� Eu���eB���إ�� ������(�s�L�^��p�������9�	anonymous�� ����e�w��� t�������� =�(:L^��� �������9K ]6/qZ/�~/�/�/ �/q/�/�/? ?C/ D?�h?z?�?�?�?� //1/3?Og/@ORO dOvO�O�/�O�O�O�O �OOQ?_<_N_`_r_ �?�?�?�?�__)Oo o&o8oJo�Ono�o�o �o�o�__%_�o" 4F�_�_�_��o� �_�����o�B� T�f�x�����o��ҏ ����Sew��� t��������Ο��+� ��(�:�L�o���f��������ʯ?Ώ�EN�T 1e��� G P!a����	� F�5�j�-���Q���u� ������Ͽ0��T� �x�;Ϝ�_�q��ϕ� �Ϲ����>���t� 7ߘ�[߼���ߣ��� ��:���^�!��E� ��i����� ���$� ��H��l�/�A���e����������QUI�CC0����!1�72.26.29'.891G#���	2�s���!ROUTER���!7`���PCJOG7�!192.16?8.0.10?CAMPRT�c�5 x1���RT� ��%/�NAM�E !��!K�JLTVL411�630R01RS�--KU1�S_�CFG 1d��� �Au�to-start{ed2�FTP=��!T�V��/��?? 1?C?U?��y?�?�?�? �/�?f?�?	OO-O?O ��/�/�/�O�?�/�O �O�O __�?6_H_Z_ l_~_�O#_�_�_�_�_��_o�o 	SM<����O�_to�O�o �o�o�o�o�_( :Loo�o�������� �2�D�� ZC��og�y������� Z�ӏ���	�,�-��� Q�c�u�����THC�� ��'�I��4�F�X� j�5�������į֯�� {���0�B�T�f��� ß՟��ҿ���� �,�>�	�b�tφϘ� ����O�������(� s��������ϔ�߿�� ������ ���$�6�H� Z�l��������� ��5ߛ�Y�k�D��� [��������������� 
.Q���dv����4(_ERR� fF*��PDUSIZ  \ �^w���>W�RD ?�%:���  ba�ckup�guest�Tfx���3&SCDMN�GRP 2g�%;� �:�\ �kD?K� 	P01.05 8��  ��  �� ��]  N�w��� ����y���2; �����������+-(�  3��v@<+/=&�9���V�����? �S/�  �
�  �s#�� �{/�j����(���S�#�� U�/� 5Vn 9S`��d/�!/�/E/2���1?234567&�? ��?�?�?O�?*OO NO9O^O�OoO�O#;�O �O�O�Oy?�?�?F_�O V_|_g_�_�_�_�_�_ �_o�_	oBo�Ofo%o �o__)_;_�o{o �o,)bM�q ���Io���(���_GROU�h*�	-0�	�!�1�cz���B�QU#PD?06��C����TYv �� T�TP_AUTH �1i� <!iPendan�������!KAREL:*$�-�?��KCT�d�v�L��VISION SCETM�ԟ��\J� �ٟ�I�'��?�9����]�o��������C?TRL j����
 .{?FFF9E3ȯ8��FRS:DEF�AULT2�F�ANUC Web Server2�
�,>۬����Ŀ�ֿ����WR_C�ONFIG k�� f2��IB�GN_CFG il��2\ @\ o<#�
~�BH|�C��?4:�~�L�DEV�`��V�>� IO ma�I��EXDAT n|����EXFLG����T�FIL o�����O�TP p�YݮaR!B���R ����	MERCA�TOR!RECO��� "R_ACHS^��ISTW*�V��,�V� "SENS�P��TXQ��990 	K�eine 0�k �h�\%IBSaC����M�4�8�@�EW�𛩀�T�L_MTN  ���� ����������l�X�SBAD��� 7�^�x�T�DL_CPU_kPCQ�\B�B���� AL��[�M�INd� =D-�T�GN��O�H����рINPT_S_IM_DO������TPMODNT�OL�� ��_PR�TY����Q�OLN/K 1q�@9�K]o���M�ASTE����SLAVE r����OZ���UOxv �CYCLu��$�K�_ASG 1sY������aП՗�~���`�$0c�������a�� ����%/0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b?pt?�?�XNUM��z��IPCH?���O_RTRY_CCNQ�I�D�N؁��8�� �Zt��FO�T�S;DT��OLC������$J23_DSP_ENB�0��ь@OBPROqC�C���	JOGI��1ukL�ad8��?����O�??"�ۯ4_�pQJ_o_ �_�_R_�_�_�_�_�zO�y8!�O-oo )_;_�_�o�o�o�o�o��o&oJ�B1 +oeNaoso�o�� ���(�:�L�^�9���BAc������ ���*�<���`�r� ����q����C����?��BPOSF�OF�K_ANJI_� K��&�RE_�.Av/���/�����KCL_�L��2�?�EYL_OGGIN7��������$LA�NGUAGE �����ENGL�ISH ١�LG�-Bw �S���S�xJ ����B����S��'� ���Z��MC:\RSCH\00\Xﶠ��?ISP x���0��⍊�ߡOC��j��Dz���AݣOGBOOK yY�$�챟X x�	��!�]�x���``͛ѧ��ه	ε���>��ϼ̲_B�UFF 1z(A�ϟ��ߞ /� �K�]ߊ߁ߓ��߷� ��������,�#�5�G��Y��}�����DC�S |ؽ =��͑�L���$�6��H�Z���IO 1}"cJO�������� ����������#3 EWk{���� ���/Cn��ER_ITMhNd ��������/ /,/>/P/b/t/�/�/ �/�/�/�/�/?��q�SEV@�mTYPhN�l?~?�?=��RS�0����B�FL 1~|�@��OO(O:OLO^OLpO�?TP��y[2}��NGNAM]���6ˢ��UPSc�G�I�0c����A_�LOADPROG� %�%UP�023}O��MAXUALRM�ܑ���筥
DR�A_P�R�Dܐ³ڑDPCf�ع�ͪ_$�;Y��P_GRP 2���[ �S�2S�	�[1�ڐ+  ��_���R#oo oYo K�Go�oso�o�o�o�o �o�o*<`K �gy����� ��8�#�\�?�Q��� }�����ڏ�Ϗ��� 4��)�j�U���y��� ğ���ӟ���B� -�f�Q���������� �ǯٯ��>�)�b� t�W������������ ݿ��:�L�/�p�[����=WD_LDXD�ISA�@+;l�ME�MO_AP�@E {?�K
 T ������&�8�J�\��n�DPISC 1��M��ϻ��T�Q���� �����2��V�h��� w�K���������
� �����R�d�O���o� ��-���������*���C_MSTR ��,=ISCD 1��͠�� ����:% ^I�m���� � /�$//H/3/l/ W/i/�/�/�/�/�/�/ ?�/?D?/?h?S?�? w?�?�?�?�?�?
O�? .OORO=OvOaO�O�O �O�O�O�O�O__<_ '_9_r_]_�_�_�_�_ �_�_�_o�_8o#o\o�Go�oko�o:MKC_FG �X�o~gLTARM_�b݅X�b ��c�� (t�b_G�RP_DO ��X�a����L��uq>k�����o$MM�ETPU��Xs���`	NDSP_CM�NT��`�Q  �I��q�al�v��_POSCF"��fΉ�RPM!���ST�OL 1�X {4@�`<#�
�� �a�� �����"� d�F�X���|���П�� ğ����<��0�r��\��SING_C�HK  %�$M/ODAQ�c��o>��i��DEV }	X
	MC:C>��HSIZE�͚`�Ȭ�TASK �%X
%$1234?56789 M�_����TRIG 1�
��lX%�ܪ��c�� Կ����˿Ͽ�<�� ��7τ�+Ϩϋ�aϣ���ϗ������/�YP����`��EM_�INF 1�w� `)�AT&FV0E0�%ߜ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����D���AL�t�/������ ����߸� ����M� �q������ Z���������%�� ��[� �2����h� �����3�W >{�@�dv� �/�//f@/e/ �/D/�/�/�/�/�� ?���a?s?&/�? �/�?v?�/�?�?O�? 9OKO�/oO"?4?F?X? �O|?�O�O6O#_�?G_�_X_}_d_�_�nON�ITOR=�G ?���   	EOXEC1�c�R2�X3�X4�X5�Xp��VU7�X8�X9�c�R kBOd�ROd�ROdbOd bOdbOd%bOd1bOdP=bOdIbOc2Vh2bhU2nh2zh2�h2�hU2�h2�h2�h2�h�3Vh3bh3�R��R�_GRP_SV �1�q� (d������5r?��>Vvտ�FN?͇��Ze�B���~e���0���U7�_D@R����PL_NAME� !>�Y��!�Default� Persona�lity (from FD) �T�RR2hq 1����Y�  	 d� ��ŏ׏�����1� C�U�g�y���������@ӟ���	��+�2�� K�]�o���������ɯۯ��<:��)�;� M�_�q���������˿�ݿ�   ��\  �  ���  ��  �A�  B�T*���
��
��@?��  �����B�p��  �C�C�P �Dz  E;� E@ D��c�C�J�q�X��d�Y�@p�t�l�`�u�e����0��d�\�]�E/~ĉ�0\�����`@o�e�0�`ż� �E	נ����^Ì��t�\�@�8T�|���EZ��å��]�|�Yũь� E Y��ߧө������¡���]����ө������� /������� �D�M�a���q�]�������T�E�  ������]��/��� -�O�Y�M�s���������������� �V�A.�E]��  ��sP�>P�d�tl ~c��! �����2 � 'EKi����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?-�F?X?j?|? �?�?�?�?�?�?�?� O0OBOTOfOxO�O�O@�O�O�O�O�M3 � �O\)�_E_���c_ u_�_�_�_�_�_�_�_ oo)o;oMo_oqo�o R_�o�o�o�o�o %7I[m�� ���o���!�3� E�W�i�{�������Ï Տ�����/�9O� ]���k����!�� ����s!�C�9�g� ]�o����̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�??X�j�|ώϠϲ� ��������O�0�B� T�f�xߊߜ߮����� ����_�%_>�P�� t����������� ��(�:�L�^�p��� ��c��������  $6HZl~�� ������ 2 DVhz���� ���
//ן9�O/ ]����/���/�/ɟ۟ �/?��??'?9?W? ]?{?���/�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_?�X_j_|_�_�_�_ �_�_�_�_�S_0oBo Tofoxo�o�o�o�o�o �o�o��,7�P� t������� ��(�:�L�^�p��� ��c��ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟����� �2� D�V�h�z�������¯ ԯ���
���/9/K/ a�o/���/}����/3� �/ω?�?�?3�9�K��y�oϝϨ��$MR�R_GRP 1��������� � `� �o ������ @D�  ��?������?������@�T;g�Ũ���*�;��	l�	 �����X�'���F�O��^ �,X� �k���K���K��eK����K~o�K{GK�M�sA�S���߈��?�;g?�����@
����Р����I����
��}v=�����X����4  �p  ?�
=ô7����A��  >�L���������	�������Ѡ����(Ѵ��,  �p�  �2����������������	'� �� )�I� ��  ����:��ÈM�È=��9�e���@u�{� v���������������������@��?��@�t��@��@�)��C~6�B�  CfK �B�B��Q������CR�Ԙ� ��� *�ވ� H�B<�� �� ����Dz��O��$�J!��� �qxy�jz  ȅ�:y�� ?��ffؿ��O G���,68��@/(*	ѝ�=$0(��V%P_(z��U�UԿ��>�33��6;���;aʤ;r��@;��;�?	�<$D���/��A0�+���?���� ?fff�!?y&02A�5@�,%5iq1 �-��]?��|?�'A� ��?�?�?�?�?�?O�OAOSO>OwOhF5F� fO�ObO�ON?�O�r9�O+_�HD�� �E�J ��E9� E��,_{_f_�_�_ �_�_�_�_�_ooAo ,i��nm2o�o�O�oX��5��Ǆ-A�G�:�F^� �E���LB:�)o&8�(:��?���_s9�B�@������yA� A��t<�	� ���7��[�F���A�d�k�����1��<���k��C����`G Ca���j~��~��}�!� �5���CHf�CW�F�B�1B-v��=���%������XR��ǽu���z�����������AP���Blz��X���}�sp��R��d�
Ák�BoU(������F<�rѵ��JGp@�KÌH�� �I%K�Ab!��L�)-yL!�GK�ӕ#HP� H��R����(��L&��J�3$�H㞀H���A��|�j�U���y� ����֯�������0� �T�?�x�c������� ҿ�������>�)� b�M�_Ϙσϼϧ��� ������:�%�^�I� ��mߦߑ��ߵ��� � ��$��H�3�l�W�|� �������������2��/�h�S���w�G��E*��~�C�?�<����Ć�����CV��L7�\]G���z_�(��`����!����1V���A3>�8!3A��vM_���v3�g��y�!�;�%D93ҵ������	/�-/,�C %P�"P_.na{o�/���/�/�/�/�+� �/�/(??8<�8?G?
n`8"�ta?#?�?�? �?�?�?�/mo'OOKO9K�QO[O�OO�K�O��O�O  �e 3��O�O__�9_'_]_kZ  2 �D��E�gE��Z�B
��q
�C)��Aj@�j�Ϝ�_�_jD� CD�0ov;j�_@�_zo�o�o�oj?`T�aZ��4jj��1jyVZ�
 �o,>Pbt ���������[��a ��I̿���Ld��2NA� @D<�U�?ϐ]� � `��a�j�A�XU�Ij��;��	la�\!��ો��e��0F��a������5���'��0Ci �P������_��?����ǟ��,nP�P���V_�z&'��9�G���k����+UUp�s�=��ͭ���Y�Ϡ�Rۯ�Z�&f���G�TY3�>��u0  '  [�e�Z�B�@�A�[��� u�R��ҿb�B�P�� @�Q.�abCp!��Tϛ�x�cϜ�ćυ�j����  �j:v�a�`x#a����
�߮� �R�dۖ��0yߋ�> Ρ�P��������쿢#>Lס ���Ao���4��e�QG�a�*��?fff?-�?& g��σ��Yb��]v�]� ��[���L桄x���� 5� �Y�D�}�h�����8�����_ F�P�� ��7��X��*� &������� -Q<u`�� ����N/r;/ �_/q/�/�/4�/�/�V/�/�/?�/7?"?�R�_4�Qn�,?�?|= (�0�~?�?�?O�? O 9O$O]OHO�OlO�O�O �O�O�O�O�O#__G_ 2_k_V_h_�_�_�_�_ �_�_o�_1oCo.ogo Ro�ovo�o�o�o�o�o 	�o-Q<u` �������� �;�&�8�q�\����� ����ݏȏ����7� "�[�F��j������� ٟğ���!��E�0� i�{�f�����ï��� ү����A�,�e�P� ��t�����ѿ�ο���+�R7(�����M�_�I��mϣϑ� �ϵ�������!��E�@3�i�Wߍ�{ܶ5P%�	P����4���B� ���	�B�-�f�Q�� u����������� ,��P��߹����� ������������ B0Rxf����  2K�� *<N`r��������/"/8A�F/T*
 T/N7 �ߓ/�/�/�/�/�/�/ ?#?5?G?Y?k?��t/���{J��4�� ���1 @D��  �1?��3 �� `?7 �27 A�X�5���? ;�s	l�2��}�K�C�0"K> F���0�?/.�?:&�uO�L > �8�ObO@/�O�O_ �O%_]�0@J_XW�x_��AЙ_�X_��_U+UU�_�_=���okiS/`�09oGh�R&f]oom�2��	�o6^u0  '�o�h�_�o_x,0�2ZO2�hB Px~� @�`�u�aEC���o��o������R�p&�4�  %��r:h&Nq~U�2��|j�|�� �в�ċ�q8�pڏ�>.a�0�1�z2�$�LƂ">L7a��pA�@=���;����s�2�3|�2�p?fff?�p?&ǐ���t�2 �4�y�5��8=���D ؟q�\���������ݯ�ȯ����7���Ffp&�s�"������ 2���뿆����3�� W�B�Tύ�xϱϜ��� ������~_,���S߮� t�ҿ��߿������� ��
���O�:�s�^�l���AfpA�����������ꈕ�o ��?�*�c�N�`����� ����������); &_J�n��� ���%I4 mX������ �/�3//0/i/T/ �/x/�/�/�/�/�/? �//??S?>?w?b?�? �?�?�?�?�?�?OO =O(OaOsO^O�O�O�O �O�O�O_�O _9_$_ ]_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Voho�o�o�o�o�o�o �o1C.gR�zvw(����� �{�����'�� 7�9�K���o�����ɏP���ی�P��P�.��~O��xT�~� i�����Ɵ���՟� ���D�/�h�S���w� ��W���=��� � 6�$�Z�H�~�l��������ؿƿ��� �.�  2��T�f�xϊϜ�@�����������C� (�:�L�^�p߂ߡ�����
 �ߒ����� ��)�;�M�_�q��������������7{J������� @D�  ��?�� � `�?��!��A�X���I� ;�	l!��}�k�e�%�<����F���K�������������=� ����=(aL� p�y���������z+v�+UU03=���m����&f�����~�u0  '/ '(K/vo/��.��̒/Z(B �/�. c@[ �%[!EC0� _/?[/8?#?\?G?EqO0�?�7  �O2I:�֮!�!�W<8�?�?n? �OD$KV18O0:OHJ>���)�M:�?�O�/��>1L��V0A��O�?�O�?O3!��!�� �?fff?� ?& 'PR?C_O4.�"Q.�M9 �}_��_Va�8_�_ �_�_�_oo=o(oao`so^o�oR]`F�  �o�o�o�on_�Y�o K�ooZ�~�� �����5� �Y� D����R���ԏ2 ��n��1�C�U��Oj� |������ӟ�����[A� A���'� 0��T�?��E�>��� ��ï��������� A�,�e�P��������� ���ο��+��(� a�Lυ�pϩϔ��ϸ� �����'��K�6�o� Zߓ�~ߐ��ߴ����� ���5� �Y�k�V�� z������������� 1��U�@�y�d����� ����������? *cN`���� ���);&_ J�n����� /�%//I/4/m/X/��/�/�/�/�/�/�'(y����?;	? ??-?c?Q?�?u?�?�? �?�?�?O�?)OOMO�;Lv�P�BPN�� {��/�O8�O�O�O_ �O&__J_5_n_Y_k_ �_�_�_�_�_�_o�O y�Co��LoNo`o�o�o �o�o�o�o�o8�&\J��w  2 o������ �2�D�V�d�����������Џ�o��
 ��]OS�e�w� ��������џ������+�{B4���{J���$MSKCF�MAP  -�?� wvD��E�  ]�ONR�EL  qE�t��p]�EXCFE�NB��
r�����F�NCƯ��JOGO/VLIM��d����]d]�KEY���=�_PAN��-�\)�]�RUN���]�SFSPDT�Y�@Ȧ����SIG�N����T1MOT����]�_CE_�GRP 1�-�t�\��	��-�?� �Oc��sϙ�PϽ�t� ���Ϫ��)��M�� q߃�jߧ�^߱����� ����7���[��P����H��l�]�QZ_�EDIT��n���T�COM_CFG 1�j���)�;�}
��_ARC_â�qE�UAP_C�PL_�դNOCH�ECK ?j� pE������� ���� 2DVh�z������NO_WAIT_L�����װNUM_RSPACEg���=�7�A�$ODRDS�P^�ѨOFFS?ET_CAR�����tDIS�rPE?N_FILE����=���SPTION�_IO#�5��M_�PRG %#%�$*/".�WOR/K ����hpIG@S% �mDC�'��m ��m!�	 ���m!<�����TRG_DSBOL  -���z���/��ORIENTkTO����C����s�A rUT_S/IM_D�q�D��TVXLCT �#B�@-5_PEsXE�g6RATs0�	�ѥx�k2yUP S�<>%�.���?��?�?OI�$PA�RAM2೏����&3	 d��VOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_���_�_o#o�5oGoYoko}o�o��< �_�o�o�o�o& 8J\n��O x������  ���  ��  A��  B�p��B���3�pH�p� g ���p�pB�p�p�p� 0�!(�P �Dz  E;�� E@ D���C� 0��q�����p�������`)�+���r �E/!�`,��qc�p���@�`����_���E	��C�/���/������p��q���EZ�n��H� ���uL��� E�qX�J�L�t���;�D�p� ���n�L�c�p���� ғ����p� d������d�� ��(�:�L�L��qE� �������� ���ҧ L�Я��q��(�:��L�^�p��������� 	�o���p��3���!��D�R�ĽĽ���p�� �ǰ� �ϸ��������.�DO ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }�������_���� ��1�C�U�g�y��� ���o��������	 -?Qcu���# 1�x��0��}�<� *<N`r� ������// &/�J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?9/�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�Oi�˿ݿ �O�_%�_M_[��O Ϙ_�9���_�_�_ oo/oE�^opo�o�o �o�o�o�o�o $ 6HZl~��� ������ �2�D� V�h�z�������ԏ ���
��.�@�R�d� v������������ �?�*�<�N�`�r��� ������̯ޯ��� &�8��\�n������� ��ȿڿ����"�4� F�X�j�|�K��ϲ��� ��������0�B�T� f�xߊߜ߮����O�O ��_C_)�7_1�[_m_ �ߘ���-o������� ����Eo��p����� ���������� $ 6HZl~��� ���� 2D Vhz������ ��
//./@/R/d/ v/�/�/�����/۟�/ ��?*?<?N?`?r?�? �?�?�?�?�?�?OO &O8O?\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_KO�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o{��� �C�)7�!_m� �o��-�?�)�������A��q�$P�ARAM_GRO�UP 1�g�X���L�`8� �o ��q��� @D�  ��?������?�p���qC�>�����t�  �;�	l��	 �����X�΀π����^ �,�X ���pH����H�ffH� � H��H�WH-���|�#�o��oi���qB�  B��������������s�4  �p � �
=É�����������ȟ�sAſ8�¼r��q�'��C���r,�2����G��wρ[��|,�  � �  �������M  �Д�����u	'�� � ТI�� �  �=�l�=��������@�"����F�������[�i������������CݐB���f������б���Ŀֿ�   ���CR>���U :��<�H�wB�pL�+�Xŷ� 3�tŕqDz�������������Ȯ�� ��x ��!�  M�,�:˅�!D�? ?�ff{R�<d��� ���ߪ���8�����ڰ�D�����(����P�!�A�x����f�>�33}����;��;a���;r�@;���;�	�<$1D4�q��A0s봂���?3�q�?ff�f��?&����A{���@�,�� ��©ᵄ�ɤ���� #���脃�X�C�|�g� �������������� 0T?x�����q�mD�� E���j E9� Eԉ��"F1j U�y����� {�-�:/�[/��/���/�/�/�/{���G?��|�3��BAȀ�/=?(?a?L?�?p9A+�A�4㠰1�?;��y?�?u?O�<?�A�OOKO6OaI����k^OC����`G Ca[OH*%D�%@�$A�A@I�ܾ���CHf�CW��FB�1B-�v�=���̞������XR���u�!_DA��ę�����AP��Blz���X��$_0���R�d�
Ák��BU(�������E@K���J�Gp@KÌH��� I%K�A�	�aLL)-yL!��GKӕ#HP?� H�R��_�P�(�L&��J��3$H㞀H���A��_#_o �_5o oYoDo}oho�o �o�o�o�o�o�o
 C.Syd��� ���	���?�*� c�N���r�������� ̏���)��M�8�q� \�n�����˟���ڟ ���#�I�4�m�X��� |�����ٯį֯����3��G���b�%�C�?�c�j�Ć�y����CV�������޿�����O�:�s�^�(d��`3��{�4�����dŏ�1V�Ϯ�^�3�>��������v��߰�v3�g� �2�!�;��%D93ҵ� L�Lٌ�z߰ߞ�����.^� Pl�P�!"//��;�e�P��t���������Q�������8�0t� ��S�>�w�b���B�/0������������8&HO�HZ  �e 3�t�6���� � 2 D�7EY� 1���B�1L�1�0C��@��A���@�?z���D� D��������/!/3/E/W/��Q?�p!������)����� ��
 ^/�/�/�/�/ 	??-???Q?c?u?�?p�?�?���! ����o̿����K�:&��1 @D�0�1y?vPA � `V��By��4�1�2L;�s	lB��RK�LC@iK��F���02O�?�O����O�LF��Ci�O�O���i�&_��J_5_n_YZ, ��@�_�V��_!��A���_�Xa_o]U+�UUoo=��� Tofk cv`�0�o�hb&f�o�m�2�	�oU^u0  '��v`B��o�oo[�B�OyAxBU��|� @e�t4C �F�B�
�C�.��,b6�m�{�  �6�:�"�!� �B�>���ÏU� ������=�+� �2�> ua�0V�=�y�k��I�#>L~a�T=�A�����ۏi%	A�3B�p�?fff?�p?& �9�*�6�B	�D4� Ed�H���HD��� ��ܯǯ ��$��H� Z�E�~���g�����ؿ O�q�s�ѿ2�ͿV�A� z�eϞωϛ��Ͽ��� ����@�+��_s�9� ���������U��� *�<�۟Q�c��ߖ��P�������T�� Q_��8�#�ϕ�o%� ��q����������� ��(L7p�m ������� H3lW�{� ����/�2// V/A/z/e/w/�/�/�/ �/�/�/??@?R?=? v?a?�?�?�?�?�?�? �?OO<O'O`OKO�O oO�O�O�O�O�O_�O &__J_5_G_�_k_�_ �_�_�_�_�_o"oo Fo1ojoUo�oyo�o�o �o�o�o�o0T ?x�u����w=(�q����� �&��J�8�n�\�~� ����ȏ���ڏ���(4�"�]�P̒Pf���b�����x��ş�� �ԟ���1��U�@� R���v�����ӯ���� ��`�*���3�5�G�}� k�����ſ���׿�����C�1�g�u�  2�ϭϿ������� ��+�=�K���o� �ߓߥ߷��������
 ����D�:�L� ^�p������������ ��b����{�J�_�+�[�~H� @D�  \��?�b� � `?��h���C]�\�X���� ;�	lh�c�}������l�����F��������+����.�Є�N	�� �o����]������]�Y�.��@N�r�+UU<wz=��ʹ��`�X���a&f�/-N�[�:/�u0  '`/n(a�/���/�u��/�(By �/> @� 45�!ECw��/[?�/ ?j?�?�?��0�?.�7  Ȗ2:�S��!%h��<O#O�? .�YOkK�18�0�O�J>�I�p�`�:�?�O�/)�>L�Sĝ0A��ODO�O<OĖ3h�N�h�10?f7ff?40?&nP�? �_�4u�iQu��9d��_ b��_SV��_oo<o 'o`oKo�ooo�o�o�o �o�o�o�o8�_�_ �_1�-���� ���4��X�C�|� g�����%ӏ����U �yB���f�x����� ;_��ß]������l>�)�A0A�f��n�w�6�����/U7/ ���ѯ
����@�+� d�O���s�����п� Ϳ��*��N�9�r� ]�oϨϓ��Ϸ����� ���8�J�5�n�Yߒ� }߶ߡ���������� 4��X�C�|�g��� �����������	�B� -�?�x�c��������� ����>)b M�q����� �(L7p� m������/ �/H/3/l/W/�/{/ �/�/�/�/�/?�/2?z7($1���T? f;P?�?t?�?�?�?�? �?�?�?(OOLO:OpOP^O�O�L��P,RP�N Q¤%?�OI8�O%_ _I_4_m_X_�_|_�_ �_�_�_�_o�_3oo Wo�O���o䈓o�o�o �o�o�o%I7�Ym����w  2Ro���1�C�@U�g�y�������� Ϗ����)�HoM�[�
 [�9��O�� ����П�����*��<�N�`�r��B{���7{J�������B��� @D�  ���?�£ � `?>�Ȣ>�C�����F>� ;�	lȢ�A}���̠)�E�F����6���A��|���E�䨮�i� G��Ͽ��,�ͽ�� �Q�_ǽϹv���РϮ�!����+UyU����=���߀&���6и�@�N���&�fd�vݮ��y��=�u0  '������ �����բa�9���B W�� @����EC�A��@������������\-�;�  ���:o�$�qU��uȢ��q���� �@����"��8������>5ѩ��С��9�+S>L>ѳt��A�D��B�����Ȣ��Ȣ��?offf?��?&�  �����բ�դ��ĥ $¨D���xc ������// />/P/'/t/_/�/ 13�/�/�/??:? %?^?I?[?�??�?�? �?�? O�?��3O�?ZO �/{O�/�OO�O�O�O �O�_#_�OV_A_z_�e_�_�_Am�A��T��S�_�_�_�Z� ���_Fo1ojoUogo�o �o�o�o�o�o�o0 B-fQ�u�� �����,��P� ;�t�_�������Ώ�� �ݏ��:�%�7�p� [��������ܟǟ � ���6�!�Z�E�~�i� ������دï��� � �D�/�h�z�e����� ¿���ѿ
����@� +�d�Oψ�sϬϗ��� �������*��N�9� r�]�oߨߓ��߷��� �����8�J�5�n�Y����}�(����� ���������
���.� �>�@�R���v��������������eP�P&=A"d��V��[ �p������  K6oZ� ~�^ O�DH�� /=/+/a/O/�/s/�/ �/�/�/�/?�/'?7  2�[?m??�?��?�?�?�?�?�?J J?/OAOSOeOwO�O��O�J
 �O�G �O__0_B_T_f_x_��_�_�_�_�_"�O���{J��$PA�RAM_MENU� ?�U��  DEFPULSE�[�	WAITTM�OUT/kRCV�Bo SHEL�L_WRK.$CUR_STYL-`{nlOPTA9a��oTB�o�bCioR?_DECSN:` �l�o�o1,>P yt�������	�aSSREL_�ID  �E1���USE_PRO/G %j%�j��CCRF`*�1c�}�_HOST �!j!����w�T 7 ��ۃ����݃�>v�_TIMEDb*����`GDEBU�G(�k�GINP?_FLMSK@�o��TR~� q�PG�A�� _��I ����CH}�  ^q�TYPEl@��4�]�X�j�|� ������į����� 5�0�B�T�}�x����� ſ��ҿ����,� U�P�b�tϝϘϪϼ����q�WORD ?�		FOL�G-c	U�	�MAKRO+�SUWCHL�C2�S7�T�TRACECToL 1��Uaw
 �@\ ]�@� � �{��2�ߗߩ�S�DT �Q��U��o�D� � � ������������*�����������������������������@���������ސ��!��"��#���$��%��&��'���(��)��*��+���,��-��.��/���0��1��2��3���4��5��6��7���8��9��:��	q�A]��+1m��Pm�k�b�o�j�Ek�k�s�m�	k�
k�k���o���o����_��_��_���������	q�	
		z� ��� b��� ���Z9�A��q��y����������O R㵼Y�a��q���y�������������� ��� ���  ��� ��� ��� ��  
�� �� �� "��  *�� 2�� :�� B�� @J�� R�� Z�� ;�U<�=�>�?�@��`��`��`�'��-`�F�\��H�I�J���B��M��`�6��D���Q����S�F`�U��L#/ "#�q�? z�? ��? b� ? ��? ��? ��? �� ? ��? ��? ��? �� ? ��? ��? �? 
� ? �? �? "�? *�? 2�? :�		��	��	��� ��� ��� ���� ��� 	��	 �� 
�� �� ��  "�� *�� 2�� �%ZU�A
q����������4		�6*����r���z����5b��Ђ�I� ���Ъ��к�������L�/ �/ �/ ��/ �/ �/ �3L��4L�4L�4L�L*IL	DLDL��/ �CL��/ ��L��L���L�L	�L�L��L!�L)�L1�L�9�LA�LI�LQ�L�Y�La�Li�Lq�L�y�L��L��L��L���L��L��L��L���L��L��L��L���L��L��L��L
��L�L	�_�+$�UL!�L)�L1�L9�ULA�LI�LQ�LY� / Z/ b/ j/ r / z/ �/ �/ � / �/ �/ �/ � / �/ �/ �+O=O|OI1� :q�U:y�:��:��:��U:��:��:��:��U:��:��:��:��:���`��`
��`� �`��`"��`*��`j2�`:��`Z:I��`R��`Z��`�:i��`r� �`z��`���`���`���`���`���`���eǰ����1� �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�k���e o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� �ek����� %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o��o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�����/�A�S� e�wωϛϭϿ����� �����o=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?1�?�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y�����s?��ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� ���������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o�� 1oWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c��u��$PGTRA�CELEN  �v�  ���A`ȋ�_UP �����������y����_C�FG ���T��Aa������Ā�����������D�EFSPD ����@a��Ћ�I�N��TRL ������8��V�PE__CONFI����ş������#�LID�á��~��GRP 1��� �v��CH������AaA�  G�G� G�7�F�,� A�  D	���A`d��)�9�~��� 	 �8���S� ´��n��B����������������B>Áe�G�Y�C� <,1<49X^� ��Z�����������v�� 9��IoZ�z�����
 B��8R@Œ���(EAL�PG���*H�=�H�x�����=(Ms^  >?V��>V�%�@����/^�!���
V7.10be�ta1� @��33@2�\@�;�CRA`C C_>  CW��T#/D�� j"0�g!}���� Dj\ �2 ��B�\ S C�] �p���!d���CX(�A�> ๙�B� ����!A��ffB�33A�33����k¶����*T"���/?��C�&�8�ѩ�� [?�?j?�?�?�?�? �?�?�?!OOEO0OiO TOyO�O�O�O�O�O�O _�O/__,_e_P_�_ ܳ �_�_n_�_�_�_ oo=o(oaoLo�opo �o�o�o�o�o�./T#F@ >y:}N`|~ ?�&�� ����/�??/?A? J��on���k�����ȏ ���׏����F�1� j�U���y�����֟� ӟ���0��T�?�x� ���_����o��ϯ� �,��)�b�M���q� ����ο����1 c=�O�y���ϸ� �����	��-�?�H� �l�Wߐ�{ߍ��߱� �������2��V�h� S��w�������� ����.��R�=�v��� ����[��������� *N9r�o� �����/�a� ;Mn�ϒ������$PLID_K�NOW_M  >:%�>!�?SV �������� ��)/;/M/�q/\/n/�/�� �M_G�RP 1��� l�CR�"�g� �&�$ �0=H��@�("1 *5&?8<���	7�+a? ???�?S?e?�?�?�? 	O�?�?9O�?OuO+DV�MR�#��-T�b�C5��"�C��  ��O�N_�O���O >___$_�_H_�_�_�~_�_�_�%ST�!1W 1��"`� �0GP�^�8�R?����a�nA8�Gay�H�PKH��GP_W.k�B�8R@Œ���(EAL�P�G��*H�=�H�x����F�o  �o�o�o�o�o �o8-?Q�u@���� o�!2o)`� �C��8�J� x�n�����ӏ��ȏڏ ����"�c�F�X�j�@���������k3� (��̟-�n�Q�c��� ������������4� �)�;�M���q���Ŀ������c4�'�� ˿,�m�P�bϣφϘ� �ϼ�������3��(� :�Lߍ�p߂��ߦ߸ߔ��c5�&���<)�n6�%�7�I�c7b�t���c�8��������cMA�D  �$"c � dPARNU/M  ��"�!|��7�T_SCHN� \�
��o�����UPDo����!>b_CMP_� Q����'�S_E�R_CHK6����cO3ERS8�@��"_MOP���_��RES_�G`�� ?aC��xFB�x5Hw�Z2�����oaC�Wq(	YߋIm4H�;C��ROQV�z �����/�)/ \E���1//�/y/ �/�/�/�/�/?�/(? ?L???Q?p?6/�� Q/�?u?�?�?	O�?-O  O2OcOVO�OzO�O�O �O�O�?���?�O�O D_7_h_[_�__�_�_ �_�_�_
o�_o.o�O��\_Qo�a� no�o�o���o�o�o�����o�V �1���������^�`�^h�]�T�]���THR_INR� �S��d�d�vMA�SS� Z�wMN���sMON_QU?EUE �š���ȡ�%MJ� �2��y��4A��  @��Bʪ����	�N- U�qN�v_m�END8o����EXE�������BE��y�j�OP�TIOv��m�PR�OGRAM %��z%l�J3�k�T�ASK_IP�ߎO?CFG ����|����ODATA��1�}�@  �}���, 2 ?���ޑ��������ڑ =+ @��	R�(F�X�@j�|�����C�1��� ������ѣ��ϭ�ө� ����ڕ���&�0�(�:�.�H��:�9����  ������������ѷC��������� �y���f�Z�v�,��%���B�ٿ����ӱ ֿƶ����"�1�=�"�-۹�O�9�a� ��V�hϰϺߞ� ����������
��.��@�R�d�v�֧s�IN�FO���}�� �C
��.�@�R�d� v��������������� *<N`r��5I���� =is�~��DIT �}��@mU��C!OWER�FL��rs��RGA�DJ �}�A�  '?��3�q�m�x��U��?C�ѐ <@	�����%qq����I�J��U˒��\9fqrbb�A<t�t$&�* /" **: ""��/'#UL"G%#��!Q)Q��� q/sE/W/i/{/�/�/ �/�/�//?�/??�? �?S?e?w?�?�?�?�? �?�?�?OO+OUOOO aOsO�O�O�O�O�O�O �O__'_9_K_]_�_ �_�_�_�_$o�_�_�_ oko5oGoYo�o�o�o �o�o �o�o�o; 1CUg���� ����	��-�?� Q�c�u������f��� -��Q�<�	)u�#A� ��=�Ɵ���
// �@/ʏ܏q� ���L� ^�˯���������ܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�Dϱ�h�zό� �����������N�� .�@߭�d�v߈ߚ�� ����������*�<� N�`�r������� ������&�8�J�\� n�������������G ��"4�Xj| ����
C.l� v<�8�؟��� � �2������ >/P/b/t/�/�/�/�/ �/;?�/??(?~?L? ^?p?�?�?�?�?�?7O �? OO$ONOHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_o�_�_�_
owo .o@oRodo�o�o�o�o �o�o�os*< N`������ ����&�8�J�\� n��������#��G� ^h����R���ş� � /*/�6/��ҏg� ����B�T�~�x����� ����ү�����,� >�P�b�t��������� ο�M���(�:ϧ� ^�pςϔ��ϸ����� I� ��$�6ߣ�Z�l� ~ߐߺߴ��������� � �2�D�V�h�z�� �����������
�� ��@�R�d�v������� ����&���< N`r����  9Kb�l���.����$PRGNS�_PREF ����� �� 
�IORIT�Y  ݔ�����MPDS?PON  ݖ���#UT&�5&�ODUCT_ID' �"���OGGRP_TG�L$m&V&TOEN�T 1�i*�(!AF_INEE ��/�!tcp|�/�!ud�/~�!icm!?��Z"XY_CF�G ��+ ��)� #��?�?� ��?�?�5�?�?�? !OOOWO>O{ObO�O@�O�O�O�O�O_*Y#t3�� %�O_a_^�>���#�!/�:_�_��-%�X��A���,  ���_
oo.o)(�T����0"�PORT_NUM#�� %�_C?ARTREP& {<��SKSTAE' ��jSAVE ��i*	2600/H601���!�_'3?K 	�ox����ݓe@������
�|�JU��e_�  1���+ p �(aԈ��#������~�a_CONFIw0��Zg#�]�U�ޔ���0��jT�ȃPt22�֋���[��C�0U��$�q�2�։�a�����8��?z�˽��i{�=J���`&�xP>>�w!��Jz��lr@�s�R��9���N��D��L¬�������=������ŐGɘ�Օٖ���V��p�� R �����y���i��� ��_������_��U]� �A���Q�w��ۯ�� ���#����Y��=� ˿)�sυ�׿鿻��� ����U���9�Kߝ� �ρߓ��Ϸ������ ����c߭�G�Y��}� ���ߛ����)�s�� ���C�U���y�����~k2S_MOTI$ ;2�֋
�?����_��);M��`�5����x����Z+ =Oas���� ���y��#�&/ ./@/R/d/v/�/�/�/ �/�/�/�/:�/7? I?[?m??�?�?�?�? �?�?�?O
??EOWO iO{O�O�O�O�O�O�O �O__/_*O<Oe_w_ �_�_�_�_�_�_�_o o+o=o8_J_Jo�o�o �o�o�o�o�o' 9K]Xojo��� �����#�5�G� Y�k�fx���ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������������ )�;�M�_�q������� ����Ư���%�7� I�[�m�ϑϣϵ��� ��Կ��!�3�E�W� i�{ߍߟ߱������� �����/�A�S�e�w� ������������ ��=�O�a�s����� ����������� "�"]o���� ����#50 Bk}����� ��//1/C/>P b�/�/�/�/�/�/�/ 	??-???Q?c?^/p/ �?�?�?�?�?�?OO )O;OMO_OqOl?~?�? �O�O�O�O__%_7_ I_[_m__�_�O�O�_ �_�_�_o!o3oEoWo io{o�o�o�o�Q�Q�Q��e�i%�f�o�fELy �o  '��mx�c�S�e  8R�Q8_��>�� �_�_ �	��-�?�Q�c�u� ��������Ϗ�_�� �)�;�M�_�q����� ����˟ݟ����%� 7�I�[�m�������� ǯٯ�����
�
�E� W�i�{�������ÿտ ������*�S�e� wωϛϭϿ������� ��+�&�8�J�s߅� �ߩ߻��������� '�9�K�F�X߁��� �����������#�5� G�Y�T�f�x������ ������1CU gyt������� �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/���/�/??%? 7?I?[?m??�?�?�? �?�/�/�?O!O3OEO WOiO{O�O�O�O�O�O �?�?�O_/_A_S_e_ w_�_�_�_�_�_�_�_ �O_+o=oOoaoso�o �o�o�o�o�o�o�_ o"oK]o��� ������#� 0Y�k�}�������ŏ ׏�����1�,�>� P�y���������ӟ� ��	��-�?�Q�L�^� ��������ϯ��� �)�;�M�_�q�l�~� ����˿ݿ���%� 7�I�[�m��z����� ���������!�3�E� W�i�{ߍߟߪì�������%��������� �%���Ӡ��Տ  (�B��8�O����� �Ϯ������ �/�A�S�e�w����� ����������+ =Oas���� ������'9K ]o������ ����5/G/Y/k/ }/�/�/�/�/�/�/�/ ?//C?U?g?y?�? �?�?�?�?�?�?	OO ?(?:?cOuO�O�O�O �O�O�O�O__)_;_ 6OHOq_�_�_�_�_�_ �_�_oo%o7oIoD_ V_h_�o�o�o�o�o�o �o!3EWido vo������� �/�A�S�e�w���� ���я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o�����������ğ ����#�5�G�Y�k� }�������ſ��үҿ ��1�C�U�g�yϋ� �ϯ���������� -�?�Q�c�u߇ߙ߫� ���������� ��;� M�_�q������� ������� �I�[� m�������������� ��!�.�@�i{ ������� /A<Nw�� �����//+/ =/O/a/\n�/�/�/ �/�/�/??'?9?K? ]?o?j/|/�?�?�?�? �?�?O#O5OGOYOkO�}O�O�3�1�1�E�I%8�F�O�F���O�O�O�E�3�E  8_2_�18?_u_|�_�_� �? �?�_�_�_oo1oCo Uogoyo�o�o�o�?�_ �o�o	-?Qc u������o�o ��)�;�M�_�q��� ������ˏݏ��� %�7�I�[�m������ ��ǟٟ�����
�3� E�W�i�{�������ï կ������*�S� e�w���������ѿ� ����+�&�8�a�s� �ϗϩϻ�������� �'�9�4�F�Xρߓ� �߷����������#� 5�G�Y�T�fߏ��� ����������1�C� U�g�y�t������� ����	-?Qc u��������� );M_q� ������// %/7/I/[/m//�/�/ �/���/�/?!?3? E?W?i?{?�?�?�?�? �?�/�/OO/OAOSO eOwO�O�O�O�O�O�O �?�?O+_=_O_a_s_ �_�_�_�_�_�_�_o �O_9oKo]ooo�o�o �o�o�o�o�o�oo o0oYk}��� ������1�, >g�y���������ӏ ���	��-�?�Q�L� ^���������ϟ�� ��)�;�M�_�Z�l� ������˯ݯ��� %�7�I�[�m������������%����ʹ��� ~h��������  �"ς��8/�e�wω�� |������� �����!�3�E�W�i� {ߍߟ�r��������� ��/�A�S�e�w�� ����������� +�=�O�a�s������� ����������'9 K]o����� ������#5GY k}������ ��C/U/g/y/ �/�/�/�/�/�/�/	? ?/(/Q?c?u?�?�? �?�?�?�?�?OO)O $?6?H?qO�O�O�O�O �O�O�O__%_7_I_ DOVO_�_�_�_�_�_ �_�_o!o3oEoWoio d_v_�o�o�o�o�o�o /ASewro �o������� +�=�O�a�s������ �͏ߏ���'�9� K�]�o����������� ������#�5�G�Y� k�}�������ů��ҟ ����1�C�U�g�y� ��������ӿί�� �-�?�Q�c�uχϙ� �Ͻ�������� �)� ;�M�_�q߃ߕߧ߹� ���������� �I� [�m��������� �����!��.�W�i� {��������������� /A<�N�w� ������ +=OJ\��� ����//'/9/ K/]/o/z|r�%�)q%�&�/�&�/��/�/�%p�%  q�/?r8?�U?g?y?�  l~�?�?�?�?�?O #O5OGOYOkO}O�Ob �?�O�O�O�O__1_ C_U_g_y_�_�_�_�O �O�_�_	oo-o?oQo couo�o�o�o�o�_�_ �o);M_q �������o�o �%�7�I�[�m���� ����Ǐُ���
� 3�E�W�i�{������� ß՟������A� S�e�w���������ѯ ������&�8�a� s���������Ϳ߿� ��'�9�4�F�oρ� �ϥϷ���������� #�5�G�Y�T�fϏߡ� ������������1� C�U�g�b�tߝ���� ������	��-�?�Q� c�u����������� ��);M_q ��������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/���??/?A? S?e?w?�?�?�?�?�? �?�/�/O+O=OOOaO sO�O�O�O�O�O�O�O �?�?O9_K_]_o_�_ �_�_�_�_�_�_�_o __GoYoko}o�o�o �o�o�o�o�o1 ,o>ogy���� ���	��-�?�: Lu���������Ϗ� ���)�;�M�_�j�l�b�x���%s������N ]��͟ ��{����`���  q��b�8��E�W�i��  \�n�����˯ݯ�� �%�7�I�[�m��R� ����ǿٿ����!� 3�E�W�i�{ύϟϚ� ����������/�A� S�e�w߉ߛ߭ߨϺ� ������+�=�O�a� s����������� ��'�9�K�]�o��� ���������������� #5GYk}�� �������1 CUgy���� ���	/(Q/ c/u/�/�/�/�/�/�/ �/??)?$/6/_?q? �?�?�?�?�?�?�?O O%O7OIOD?V?O�O �O�O�O�O�O�O_!_ 3_E_W_ROdO�_�_�_ �_�_�_�_oo/oAo Soeowor_�_�o�o�o �o�o+=Oa s��o�o���� ��'�9�K�]�o��� ������ۏ���� #�5�G�Y�k�}����� ������ҏ����1� C�U�g�y��������� ӯΟ��	��-�?�Q� c�u���������Ͽ� ܯ� �)�;�M�_�q� �ϕϧϹ�������� ���7�I�[�m�ߑ� �ߵ����������!� �.�W�i�{���� ����������/�*� <�e�w����������� ����+=OZ�\�R�ht	%c��� �� � ��ttP�t  8��R�8�5|GY� L� ^�������/ /'/9/K/]/o/B�| �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�/�/ �?�?�?�?OO1OCO UOgOyO�O�O�?�?�O �O�O	__-_?_Q_c_ u_�_�_�_�_�O�O�_ oo)o;oMo_oqo�o �o�o�o�o�_�_�_ %7I[m�� �����o�o!�3� E�W�i�{�������Ï Տ������A�S� e�w���������џ� �����&�O�a�s� ��������ͯ߯�� �'�9�4�F�o����� ����ɿۿ����#� 5�G�B�T�}Ϗϡϳ� ����������1�C� U�g�b�tϝ߯����� ����	��-�?�Q�c� u�p߂߂�������� ��)�;�M�_�q��� ����������� %7I[m�� ��������!3 EWi{���� ���////A/S/ e/w/�/�/�/�/�/� ��?+?=?O?a?s? �?�?�?�?�?�?�?�/ �/'O9OKO]OoO�O�O �O�O�O�O�O�O_O OG_Y_k_}_�_�_�_ �_�_�_�_oo_,_ Uogoyo�o�o�o�o�o �o�o	-?JcLa�BaXudy%Sv}�v���t� �
��d}ds@cdu  8��Ba8�%�|7�I�� <o No��������Ϗ�� ��)�;�M�_�2ol� ������˟ݟ��� %�7�I�[�m��z��� ��ǯٯ����!�3� E�W�i�{��������� տ�����/�A�S� e�wωϛϭϨ����� ����+�=�O�a�s� �ߗߩ߻߶������ �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� �����������1C Ugy����� ��	?Qc u������� //)/$6_/q/�/ �/�/�/�/�/�/?? %?7?2/D/m??�?�? �?�?�?�?�?O!O3O EOWOR?d?�O�O�O�O �O�O�O__/_A_S_ e_`OrOr_�_�_�_�_ �_oo+o=oOoaoso �o�_�_�o�o�o�o '9K]o�� �o�o�o����#� 5�G�Y�k�}������� �������1�C� U�g�y����������� Ώ��	��-�?�Q�c� u���������ϯ�ܟ ��)�;�M�_�q��� ������˿ݿ���� �7�I�[�m�ϑϣ� �����������
�� E�W�i�{ߍߟ߱��� ��������/�:�<ш2�H�T�%C�m�w�o�ckd�� me=�T�T�0�T�  8����2�8���|'�9�� ,� >�w������������� ��+=O"�\� ������� '9K]oj| ������/#/ 5/G/Y/k/}/x��/ �/�/�/�/??1?C? U?g?y?�?�?�/�/�? �?�?	OO-O?OQOcO uO�O�O�O�?�?�?�O __)_;_M___q_�_ �_�_�_�_�O�Ooo %o7oIo[omoo�o�o �o�o�o�_�_�_!3 EWi{���� ����o/�A�S� e�w���������я� �����&�O�a�s� ��������͟ߟ�� �'�"�4�]�o����� ����ɯۯ����#� 5�G�B�T�}������� ſ׿�����1�C� U�P�b�bϝϯ����� ����	��-�?�Q�c� u�pςϫ߽������� ��)�;�M�_�q�� ~ߐߢ��������� %�7�I�[�m������ ���������!3 EWi{����� �����/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/� �'?9?K?]?o?�?�? �?�?�?�?�?�?�/? 5OGOYOkO}O�O�O�O��O�O�O�O__����$PURGE_ENBL  ,A>-A�-A4P�WF<PDO  hDT,BOQ TR_I]T�gQKUTQRUP�_DELAY ��"A"AKU,B�R_H�OT %�UiR%�+B�_�]�SNORM�AL�XKR�_!o�WS�EMI o&oeopQQ�SKIP_GRP� 1ĞUMQ? x 	 ho�o �o�o�o�o�i�U'w GYk1�}� ������1�C� U��e���y�����ӏ ������-�?�Q�� u�c���������͟����)�;��U�$R�BTIF^T�ZY�C�VTMOUT^Vv�U�Y�DCR�c}ƈi ��a�E ��E-�+�E��1C�s'�DO�DC���m�l���J� �'�������-å��2�o� ;���;aʤ;r��@;��;�?	�<$D�/@8�j�{� {��� ��ſ׿�����1� C�U�g�����vϯϚ� ������	�L�-�?߂� c�u߇ߙ߽߫����� ����)�;���_�J� ��n������ �� �V�7�I�[�m���� ���������������� 3WB{f�� ����*�/A Sew������,kRDIO_TY_PE  �[���REFPOS1� 1Ǟ[
 xSoY)�}/��/�- L/^/�/�/�/?�/A? �/e? ?b?�?6?�?Z? �?~?OO�?�? OaO LO�O O�ODO�OhO�O _�O'_�OK_�Oo_�_ _._h_�_�_�_�_o �_5o�_2okoo�o*o�oNo�o�o/%2 1�;+J/�o�oL�o pvo�/���� ���6��Z�l�-'3 1�
��V� ԏ��������@�ۏ =�v����5���Y��<p�0$4 1ʍ��� ��۟Y�D�}�����<� ů`�¯�������C��ޯg���0$5 1� ��&�`�޿ɿ�� &���J��Gπ�Ϥ��?���c���z�0$6 1�;+������`���τ��3!7 1� �.�@�z�������S8 1α��������x��/�SMA_SK 1�� H 8������XNO����4�D�/!MOT�E  �M�_CF�G �[�D�."P?L_RANGW�+!�_���OWER ��;%��g�."S�M_DRYPRG %;*%X� ��TART ����
UME_PRO�����j,$_EXE�C_ENB  <�c�GSPDC � �e��GTD�B��
RM��M�T_��T��Y��O�BOT_ISOL�C����x'N�AME ;*�KJLTVL4�11630R01�x0�O�OB_�ORD_NUM �?��
!�H6�8�895�  �+!����������|� �/ PC�_TIMEOUT��� x/ S232�t�1�;%� L�TEACH ?PENDAN�p�G�I�nW���Maintena�nce Cons�o�C�R,"b/��	�UnbenutztY*�/X/�/�/�/�/8�/�b"NPO ��K���SCH�_LF ���	��1T;MAVAI�L��5��c�SPACE1 2��
 K?HHG��v�F������4L8�?�L;WOL? ;O�O�O�O�O�G�?O O%O�OIOkO]_~_A_ �O�_�Y�#��]�O_ _%_�_I_k_]o~oAo �_�o�o�o�O�_o!o �oEogoYz=�� ���o�o/� Suw9��������� ����+�ُO�q� c�����������ߏ� ��'�՟K�m�_��� 3�������˯���� #�ѯG�i�[�|�?��� ����ǿ�����1� C�U�WϾ�;ύϮυ� �����	��-���Q� s�e�7߉ߪ߼ߓߥ��52�?�?���#��� G�i�x��\����� �����*�<�N�`�r� t���X���������� �&�8�J���n���� T������" 4F�j�~�R ����0B �f�z/�/^/��/ �/�///,/>/�/b/ �/v?�?Z?�?�?�?�? ??(?:?L?�?p?�? �?VO�O�O�O�O OO $O6OHO�OlO�O�_�O �_�_�_�_�O_ _2_ D_�_h_�_|o�oPo�_ �o�o�o
oo.o@o�o do�ox�\������3��
�.@ �d�����y�ˏ� ӏ�5�G�Y�k�}� ������u�ǟ蟿��� �1�C�U�g������ ��q�ï���ͯ�-� ?�Q�c���������� o����ٿ�)�;�M� _�σ����ϸ�{�ݿ �����%�7�I�[�	� ϡϓߴ�w������� ��!�3�E�W�i��� �߱�s��������� /�A�S�e������ �����������+�=� O�a�������m ����'9K] ����y���/�4�'�9K ]/���/�/�/�/ 	?�/?#R/d/v/�/ �/�/�??�?�?O�? O<?N?`?r?�?2O�? �?�O�O�O__�O8O JO\OnO�O._�O�O�_ _�_�_o�_$oF_X_ j_|_*o�_�_�o�o�o �_�o BoTofoxo &�o�o����� ��>Pbt�4� �������ڏ� :�L�^�p���0���ȏ ���ޟ�����6�H� Z�l�~�,���ğ��ׯ �������"�D�V�h� z�(�������ӿ���P	���#+52.D/ V�h�z�(Ϟ�������@���&��;�#+6O� a�sυϗ�E߻����߀���"�C�*�X�#+7 l�~ߐߢߴ�b����� 	�*���?�`�G�u�#+8���������� �&G
\}d��#+G �5+� �:
�   �,:5%K] o��������o�>d �%/7/I/ <j/|/�/�/��� �*�/�+?
/;?M?_? q?d/�?�?�?�/�/�/ �/?O7O*?[OmOO �O�?�O�O�O�?�?�?�O$O6_ `� @> oU�}_�O�_ �Ek_9_�_-Oo�_�_ �_�_loo1oSo�ogo �A�a�E�c�o�o! �e�oSe�9k ����������L
�_n�@�_MO�DE  ���S ��]�_ZA���_�9�	4��]�D�CWORK_{AD���c�F�/R  ����b���_INTVA�L�������R_O�PTION̖ ���F�TCF� ې����?��7���V�_DATA_GR�P 2��H�DU@PJ�y�F�����G� ʯ���ܯ� �6�$� F�H�Z���~�����ؿ ƿ����2� �V�D� z�hϞόϮϰ����� ���
�@�.�d�R�t� �߈߾߬�������� ��*�`�N��r�� ����������&�� J�8�n�\�~������� ��������4"D jX��Be����� ���q�5#YG }k������ �//C/1/O/U/g/ �/�/�/�/�/�/	?�/ ??-?c?Q?�?u?�? �?�?�?�?O�?)OO MO;OqO_O�O�O�O�O �O�O�O___%_7_ m_[_�__�_�_�_�_ �_�_�_3o!oWoEo{o io�o�o�o�o��o�  ��o�oAwe� �������� =�+�a�O���s����� ��ߏ͏��'��3� 9�K���o�����ɟ�� �۟�����G�5�k� Y���}��������ׯ ���1��U�C�e�g� y�����ӿ������ 	��Q�?�u�cϙχ� �ϫ���������o>� b�M�ߕ�߹ߧ� ���������%�[� I��m������� ����!��E�3�i�W� y�{����������� ��/eS�w �������+ O=sa�� ����//9/'/ I/K/]/�/�/�/�/�/ �/�/�/�/5?#?Y?+���$SAF_DO�_PULS  �-��������1t0CAN_T'IME�0}��3����1R �����8		��U��
�8���4�4�� ^�OO 0OBOTOfO�?�O�O�Op�O�O�O�G�1  B2T�1�1QdXQ Q�4}��1�� @CVT[�0@P_z_�\�1�_�WP�U�� @B�3T i_�_�_o~iT D��o AoSoeowo�o�o�o�o �o�o�o+=OpaX^?VNVpy 
�qp��yz�3�1;�o}���4p{}
�t� �Di�0�A�1�z?�� �B�1�q�1�A�1z�Y�k�p}�������  �������� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я�����$��h_H�Z�l� ~�������ƿؿ'�>T�Q���R�7�I� [�m�ϑϣ�Žρ�A0�22�@U<�}���@�$�6�H�Z߁�^�^ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ���������, >Pbt���#�� ���(:Ll�2��P�i%mih��0�A �B Ѓ����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO0*O<ONOYG�=X�� *`YO�O�O�O�O�O�O __&_8_J_\_n_�_P�_�_�_�Z�B��_��V�_i��A���_/m	1234�5678�r`!�B  �/h�@��jo|o�o�o�o �o�o�o�o q�O#5 GYk}���� �����1�C�T� w���������я� ����+�=�O�a�s�8����V�BH��П �����*�<�N�`� r���������̯ޯ�[�;�j��&�8� J�\�n���������ȿ ڿ����"�4�F�]�D�_wωϛϭϿ��� ������+�=�O�a� s߅ߗ�Z��������� ��'�9�K�]�o�� ������������ #�5�G�Y�k�}����� ����������1 C�gy���� ���	-?Q cu���Ug`����`�//%(�"C��A�_J  W �mH2qBgbj%)
�Pdq#�?`��R2��/�/�/�/��+pM$ZO�� �/0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O?�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ ooG!�$SC�R_GRP 1����� �t �G!� R%	 /Ra�Zbkb dd�f%f!�ekwg�o8�o�o(-�a �b?D�` D��.qc�w�k<R-2�000iB/21�0F 56789�0� @tX� R�B21 OpC#
V06.10 zpB�hKa�br#�u�vZa�fIa�cIa3f!"�ahj�a�y	�r��
��.�@�P��G�H��r�r^g�v�O	q��a4��)7'D�o��C��B������va´ �����A����A?���� �B���P�  �>����d���)/�D�mhZ`�OG!�o��o1��.'"��h�p�X��ŚeB���/B�  ~�ǐ�va9AL ��  @G ���va@�`ʟ  ?����v�: 򟨛vaF@ F�`�%�� I�4�m�X�}�����ǯ ��믖i��������%�7�B�E�گ�� v�����ӿ��п	��� -��Q�<�u��/���c�o����i
����C#�@㑬�;��hΟ�@�B�P�1234Ns`׀h���C$�A�gRa��㏛cd!2�rG! ��������2�>�P�� Pv�(|���� Ibp`�tZ` �}�{yi��gϩo�i7р�P�����7u�Indepe��nt Axes Qs	����n�f�w� �s�w3i��r���j |����c��	�v���/A�� Z��~iϢ�S�� /������/���F/ 藦�t/��/��/�/ �/�/?�/?=?(?a? P�:�p?�?�?Z��?R? O�?'OOKO6OoOZO lO�O�O�O�O�O���� #_f�����k_}_�_.�Rٺ_\�n�~�o�� L$o7o��boto�oUo �o�o�o�o�o��S�����_�� :��._��������� ������p�$6H Zߏ���'��� �o�~������Hoh ퟀ��#��G��h� 
/��./P/R/d/�� �0�1��U�@�e��� v�����ӿ�?�?��� ��?Q�Ŀu�`ϙτ� �Ϩ���������;� &�_�
�_m��F_X_ �����_�_�_�_�V�_w�o������o �������+�=��a�s���$6xBT�� ��3��W� ��,�>�P�b���� ������ΏSew� �:�L�^����// +/��ܟa/��/�/6� �/Z��/~� ?��įƯ دZ?|/�?�/�?�?�? �?�?�?�?#OOGO6�  �VOhOzO@��O8O�O �O_�O1__A_g_R_ �_v_�_�_�_~���_ L����Qocouo�2�8�J�8ff��o��4/ Z�Wi8y���������$�SEL_DEFA�ULT  ��_��P��MIPOWERFOL  6e.�7�oWFDO#� .���RVENT 1O����,��`�L!DUM_E�IP����j!?AF_INE"�Ə��T!FT����伏�!�>� ���e�!RPC_OMAINf�H��T����x�VIS��G�������!TP�P�U����d�I�!
�PMON_PROXYJ���e8�����c���f���!R?DM_SRV⯯�9gЯ-�!RZ�I����h�y�!
z�M䬯��ih�ſ!R�LSYNCƿ��8���!ROS̛�8��4 �]�!
�CE�MTCOMd^ϲ�kLϩ�!	r�OCONS�ϱ�l�� ��,�������B�g� .ߋ�R߯�v��ߚ��߀������?����R�VICE_KL �?%�� (%SVCPRG1r�D���2����3��D���4
����52�D7���6Z�_���7��D����8������9������D������' ����O����w��$� ���L����t���� ������?����g �����=���e ���/��//�� �W/��/��-�/ ��U�/��}�/�� w������B?�?�� �?�?�?�?�?�?�?O O?OQO<OuO`O�O�O �O�O�O�O�O__;_ &___J_�_n_�_�_�_ �_�_o�_%ooIo4o [oojo�o�o�o�o�o �o!E0iT �x�������M:_DEV ~���MC:�����%�~�L S  ���i��!��OUT�`�:�!�R�EC 1�d5L���   �S 	�  � � � ��ą��� ��ӎ	 �����އ��;�K5
 �W7Q6 ����`�l�d5����	M�U ��M��+ ��>��7�] �@7�������7�I �r�����������Ks�]��Y�]�XG�m��� R �� �
̑�����џ��͟�c��>�\� U�����	��Ư-� �M��P��
�� �}�g�y����$��7���� W ��T��F]��`� ��� ���� �H�Q�"M�ӯ  �M�&)��U` �?7����7��H �t���z��������
��ݢ�����υ���U� �� �m�? ��Pտ�� �sY��n�����h  -��6���]�s�T-Ϸ���' �� ���]� "��k�ѿ���a��7��!�  ������P�k�$�6�|M�� �Y� �P�� �-ߨ�)ߋ�b�'7�����T�E����X�k����m Y��L�P �dM��u��=��S� � � �f �k����M��7��7�7�KZM��5�	~ �l�oV���P�������P�e�����*B�@�� �����p��������֛��M��7�����	�����������b>�A���H�)�B�����+�����K�7���D�50�� �U��-��B� TϾ�xϊϜ���*� <�N�`�r����b� t�>�ߪ�t������ �Ͼ����������|<�N��V�� �!��C/K4�m�� ��� �V�/�� �!7��7�eG7��E��/	��o�����E��vQ�c�u�������}/�/����u��2d�/����Ā�?������2��B�@Դ]��	�0���6K^b�,�M�L�.����@ 
IO ���4D��O��  a>�D�!�?���7�~@�g���U�����,�!,��_�41�� 8 VE_ ��M�� �J �~�GOT)?;2J�_	81���� 0
��@��6�OUi�<!,��$�� � ���_ j� ��^����T�_�27��7��7�٢�uo�j� �����x��I������o"��o��� ,aT�Lb���6 ���-Mi��'��  �) ���	��SNh�`6��/�����k�����m�s�]���N�)�}{)��������S����	�g�я!��i�G�Y�ß�S"Q�ş˟���R/H"�a���o��S��q�w�a���RRk�k}p*)G'��������S�A��<e��ST�l�! �0�S�m�K�]�ǿ���ɿϿ����� %�K�9�o�]ϓρϷ� �ϫ��������!�G� 5�k�M�_ߡߏ��߳� ��������!vp�/�0��G�}�O%$ׁ�� q���)�;����)��� M��q���������`��������%��y �k����k�3
�A���-?���17!W7O�%M�_���T�����+/W7N�@=�///S/e/�2�/ �/y/�/	�/�/�/1?�?U?C?y?3�����e�?c?�/�?A�A(�?�?�?/O�0ƅ� #OOSO�O�EH��O |O�O0�L_H)__ M_8_q_�_vpe?�O�O �_�_�_o�_%o7oo [oIoomo�o�o�o�o �o�o�o3!WE {�o����� ��/��#�e�S��� w�����я�ŏ��� ��+�a�O�����y� ����ߟ͟���9� �]�K�m��������� ۯ�ϯ���5�#�Y� G�i���q�������� ׿���1��L�_,�v� dϚψϾϬ������� ��$�*�<�r�`ߖ� xߊ��ߺ�������  �J�,�n�\�~��� ���������"��F� 4�j�X�z��������� ������BT6 xf������ �P>tb �������/ //L/./@/�/p/�/ �/�/�/�/D�n_'?? K?6?o?Z?�?�_X��/  ?�?�?�? OODOVO 8OzOhO�O�O�O�O�O �O�O�O.__R_@_v_ d_�_�_�_�_�_�_�_ �_*ooNo0oBo�oro �o�o�o�o�o�o& 68J�n�� �����"��2� X�:�d�j�|�����֏ ď����0��T�B� `�f�x���������ҟ ���,��P�Fϸ?^� `��������ί�� ��:�(�^�L�n�p��� �������ܿ� �6� $�Z�l�Nϐ�~ϜϢ� ����������D�2� h�Vߌ�zߘ��ߤ��� ������
�@�.�d�v� X����������� ���$�*�<�r�`��� ������������  &8nP~�������f��$�SERV_RV [1�i���0(	 \�n���!�3TOP10 1��=
 6}�q�6 q�U �q� q�� 2q�6 �q�6 *!��?YPE  q���Hq�1HE�LL_CFG ��t&�0�? ��?�/q�%RSR �/�/�/??:?%?^? I?�?m??�?�?�?�?� O�?$O5MDD<I�
 �E%5OvO�OCE�?M2!�O�B�@�D\D1!d�Oq��)}}&HK 1�+ �O<_7_I_[_ �__�_�_�_�_�_�_ oo!o3o\oWoio{o�C}&OMM ���/�o|"FTOV_�ENBi$Et*OW_REG_UI�o~{"IMWAIT�b��I{OUTv�DyTIMu���WVAL,s_UNIT�c�vt%Q�LCpTRYw�t%1MB_HD�DN 2�k )P����� >�5�G�t�k�}������̌�qON_ALI_AS ?e�iLhep���(�:�L� D��w�������X�џ �����ğ=�O�a� s���0�����ͯ߯� ���'�9�K���\��� ������b�ۿ���� #�οG�Y�k�}Ϗ�:� ���������Ϧ��1� C�U� �yߋߝ߯��� l�����	��-���Q� c�u���D������ ����)�;�M�_�
� ����������v��� %7��[m� �N�����! 3EWi��� ����////A/ �e/w/�/�/F/�/�/ �/�/?�/+?=?O?a? s??�?�?�?�?�?�? OO'O9OKO�?oO�O �O�OPO�O�O�O�O_ �O5_G_Y_k_}_(_�_ �_�_�_�_�_oo1o Co�_Toyo�o�o�oZo �o�o�o	�o?Q cu�2���� ���)�;�M��q� ��������d�ݏ����%�Ѓ�$SMO�N_DEFPRO ���N�� *SYSTEM*Ё��>�RECAL�L ?}N� ( �}׏����ԟ��� ���/�A�S� e�w�
�������ѯ� �����+�=�O�a�s� �������Ϳ߿񿄿 �'�9�K�]�o�ϓ� �Ϸ������π��#� 5�G�Y�k��Ϗߡ߳� ������|����1�C� U�g�y�������� ������-�?�Q�c� u�������������� ��);M_q ������� %7I[m �� ����~/!/3/ E/W/i/�z/�/�/�/ �/�/�/�/?/?A?S? e?w?
?�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O�O _'_9_K_]_o__�_ �_�_�_�_�_�_o#o 5oGoYoko�_�o�o�o �o�o�o|o�o1C Ugy���� ����-�?�Q�c� u��������Ϗ�� ���)�;�M�_�q�� ������˟ݟ�� %�7�I�[�m� ����� ��ǯٯ�~��!�3� E�W�i���z�����ÿ տ������/�A�S� e�w�
ϛϭϿ����� �ψ��+�=�O�a�s����$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1z� �?��%����<�Q�����_*_�G�ֶo1�6�w� �.�f���֦����� ׯ�q#����� ���7��$�E&�g����KV���֟q8����֡0������!�0��'�� t�W��8� �� �v���/����vc��
�2�G
̈́6w��q��� ׆���� �lG�/��q���6/ �Q�&/g/�Q<V/�/�#����/h	�/�/� ��/&? ׄ���?W?I�F?�?�&�v?�?�2�Y8�?�?��ϴ�?O��׋OGO��1�6OwO��?�O�Y�|x�O�O�	q�O_�n�M�O7_��	�&_g_���߅/�_ �J�\�_�_��5O�_ �c�u?&o��5Oo�Wo�O�Eo�o �]co�vo�o�獦o��o�zb�� ��1�%/F יC�Ov�����f�:� ���7�/� ��c���7��'AJ&��g�ֵ��� ע��%��ǏւA/8������4��'���~j�W��@q��� ��I�v������>w���ZwN1�֟��R�u�F�� ����6�w��'�qf���֑�����ׯ��6�O� א��6��I|&�g� ׁ'���ߋ�̿Ѹ#����� ��'�p���]���#tF�̇�և��R��PA�RAM ����� �	�P�<�P!�I�D���OF�T_KB_CFG�  ]��ԉ�OP�IN_SIM  ����=�O�a�Q ���RVQSTP_DSB&����h���SR �)�� � & FO�LGE125 .<����0001A������THI_CHA�NGE  �E���GRPNU�M� �OP_?ON_ERR��~I�PTN )վ�C�R?ING_PR1�U����VDT+� 1	�ɑ@�@���F�� ������� �1�C�U� g�y������������� ��	-?Qcu ������� );M_r�� �����//%/ 8/I/[/m//�/�/�/ �/�/�/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O�O __+_=_P_a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o�o#5 GYk}���� �����1�C�U� h�y���������ӏ� ��	��.�?�Q�c�u������e�VPRG_�COUNT��8|��ƒENB�����M�4���UPD �1���T  
 ����B�T�f������� ��ׯү�����,� >�g�b�t��������� ο�����?�:�L� ^χςϔϦ������� ����$�6�_�Z�l� ~ߧߢߴ��������� �7�2�D�V��z�� �����������
�� .�W�R�d�v������� ��������/*< Nwr����� �&OJ\ n����������_CTRL_NKUMГ!�!"wGUN%" 2�0��  1$4!!
4!/s$
1$Ւ(#��'�/�/�/�/ÐY?SDEBUGА1��� d�� SP_�PASSЕB?~;LOG �0��� J1��^��k$[=�%?UD1:\04.�12_MPC6? (c(�?g=x82�?�2?SAV �9=�!ln%&x8SV�;�TEM_TIME� 1�R+ ( w?Z�"0����  ��>hF�qsH�O�O�O�O�O��/T1SVG S+�ѕ�'��PASK_OPTIONА�0��ߑ'Q_DI�0�ߔTBCCFOG �R+�=�.�_`�_���!�_ �_�_o�_5o oYoDo }oho�o�o�o�o�o�o �o
C.@yd ������	��%�6��i�{�� X�����Տ�����0� �=P�!�G�5�k�Y� ��}�����ßşן� ��1��U�C�y�g��� ����ӯ������	� +�-�?�u�[�F����� ��˿ݿ[����7� %�[�m��Mϣϑ��� �����������E�3� i�Wߍ�{߱ߟ����� �����/��S�A�c� e�w�������� �+�=���a�O�q��� ������������' K9[]o�� �����!G 5kY�}��� ��/�1/��I/[/ y/�/�//�/�/�/�/ �/?-????c?Q?�? u?�?�?�?�?�?O�? )OOMO;OqO_O�O�O �O�O�O�O�O__#_ %_7_m_[_�_G/�_�_ �_�_�_{_!oo1oWo Eo{o�o�omo�o�o�o �o�o/eS �w������ �+��O�=�s�a��� ����͏���_	�� 9�K�]�ۏ��o����� ��۟���͟#��G� 5�k�Y�{�}���ů�� �ׯ���1��A�g� U���y�����ӿ��� ���-��Q��i�{� �ϫϽ�;�������� �;�M�_�-߃�qߧ� ���߹�������%�� I�7�m�[������ ���������3�!�C� E�W���{���g����� ����A/Qw�e��� �$TB�CSG_GRP �2����  �  
? ?�͐��8��  <N 8r\���� ����/,//P/ :/t/�/l/�/�/�/�/ �/?�/(?:?$?^?D? n?�?~?�?�?�?�?�?�O�?6OHMA��*SYSTEM*� �V8.2306 �qC4/2x@014� A t  �_F_GF�� PAR�AM_T   ��$MC_M�AX_TRQ���$�D_MGN�CC�� AV�ISTAL��IBRK�INOL�D�FSHORTMO_LIM	Z�M�E�JPTPL1CU2�CU3CU4CU5CU6�CU7CU8�A ���A��A� ��_ACCEJRx�WTQ�SPATH�W��Q�S�Q_RATI�O�B�S�@ 2 � 	$CNT_S�CALE	ZSCL��CIN�Q_UCA���bCAT_U�M%hYC_ID g	*cB`_EKP�GjTPGj]PG`PAY�LOAWJ2L_UPR_ANG�f�LW�k�a�i�a�ER�_F2LSHRT�gLO�da�g)c�g~)cACRL_Shppgzd�BHVA`?  $H�B:roFLEX7s̝@�Jb�@ :]$aLENKQguTQ$DEjx�t|s�R�X�p�zSLOW�_AXIq$FU1aI�s2�x1�q��u�wMOVE_T�IMd_INERsTI%`:p	$D	�?TORQUE�Q!��p�IHPACEMAN�`��P�s�E^��V�p�A/�x�@�x�TCV���@��A�������@T.��@��!J�A����M	�(a|�(`J_MODa��p� R�@�Jgq2�@P�^�Eo�H0`J��Xp�A�R�U�?�JK.�����K�KSVKTSVK]SJ�J0�KSJJTSJmJ]SAAKSAATS3AA
�fSAAoS�AN1ǌ<����@�@P�E_NUQl�VqCFG�A �� $GROUP��@SK&cB_CO�NFLIC�dB_REQUIRE.q��qBU sUPDAeT�v� �ELk��� Τ��$TJ��P�JE�@CTYRa�qTN	�F˦���HAND_VB�8rVqOP�U �$]�F2�F
�TSC�OMP_SW&a�r��@�F� '$$M�`�IR�C|���A��x��R��A_�}b�FDļ�MA�LA��LA�KA [Ұ�KD��LD�KD [P�PGR�Gp�ST�Gp��IZp�NXDY�`R�@ �E��ڵ�` `�g�q�g �a�g0�<Q@��p��UPKUTU]UfUoUxU�Ur�R�Us�T r�Wt�R %�n�TPy�OASYM�U:p� ��V�Pm�ao_SHo�g4d]��C�>oPoboto�cJ�l>P�jp^�T�i
�_VI&����Ѫ�V_UN!I�c��TS�aJ���� ����l���e����m��y>P1a����GtOs ��TC�PPIR�A  >��ENABL�p�����$TCDEL�AY�R��SP�EE4P  X ��I�N� ސ��� GP����Q���q��@MPڢPROG9_���YPEڡ��_z�	 |�m���SE s��m���' Ǧ�WARNI��EN&���OTF�qj��3_T���MAARSuCW���SPDz��
 ������EA�RTBE���ET芠z���PPARGAT��FLG�u�|sUS�@E�@R&��6�%�aos6RE�AJVXTR ԱO;UT�A p렜��� E�̢�ID`�(d^�Uc�A� `��޵�G�Q# �PH���<��{�I�$DO�  s���z� �
�I��A��J �p0��W#�۠���q�� � T�M�ES���R���T� P��"@Pl� ��#��(�!�)T"�m�� $DUMM�Y1]Q$PS_f�pRF�pg@$�&��FLA|��2>�GLB_Tu�k*5���(���8!e�����QSTT���SBR�PM2�1_V�T$SV_ER�`O�p3�3CLD0p2A^�����GL��EW�A �4��$��$ZBݲW�3���`P�As �%b  `�3U�5� ]�N�0�$�GI�}$�1 ���3�0�A� L��F�}$FJ�EFN� M�NcyF]IJ�TANCb_  ��J RǱ� + $JOgINT���$�3IM� �Q��FECE�q��S�b,�*B���Q_� �pUS��?��LOCK_�FO�`[�� BGL�V��GLXT  _sXM`�AEMP�@��� -PB2�@$US�!�0p2*��4QQ�RW��@QQ�SCqEj�CrP $K���M#TPDRA8�0�T�AVEClp�V֊@IUQQVQHE��@TOOL�s�SVv�tRE�PIS3|sr�T64�)`ACH� ����QON��$2�9�"�PI�  �@$RAIL_B�OXE���RO�BO"T?�r1HO�Wc>d� aROLM�"ge_�
dxb��/`��p6�O_F��!�   �2�Q^q��O<�R�PO]r�b�p�A�` �$�3~X2MU�֡X���@	 IP#VNK���R/b�Q
�QQ�`�PCORDED�@���`��a��OY   7D )0OB�٣ �@dwSq�#E Sr�ۡwSYSSqADR �=QTCH�� S , �A�A_D��th�)"��VW�VA�� � ��P�2kPREV_�RT��$EDI}T�VSHWR�����$�K��IND�� `;�$��D�&�[�U�6��KEp��� �l�JMPpp�Lj|�TRACUE)[p�I,P5SڢC �NE�Pۡ���TICK�S��MnOF<��HNR1� @]p��L	_qGK&f��STY�vaLOD1 �@�����~� t 
�
 G�u%$�qD=:� SFp!$��8�!�F �P��LS3QUaLO����TERC� ݱ0�;TSz�:�g1@�� p��㡼Q,�O� ��#dIZ4A���! C�"!�oUTsPU��1�_DObBֿpXS�@KjAXiIP��cVQUR���0i#$TH`�~vK����_�P�rET��P( Rlp��O�F��P�A�����$ cc�>   # SR3� l:�u��a ������������ ù�ӹR���R��R� �d�~�B�d����҂�	C翐�C��� �2�D�'�ĐSC,0 o! h�0DS�4� X}�AT��<��� ~���"ADDR�ES�SB�SHIyF�HP_2CH� �zqIK0���TX_SCREEUr"	 =k�TINA�3@���D  ��`Q9_��T0# T���0 '�g00�^��r^�>�RROR_vA���(�h$ \�UE�5$$ ��Щq0S��1�qRSM��T�U�NEX��j���S_�3��G�ѽ���G�⒡C�B��� 1g# 
z��%="X�2��MT!�Lv��m�w0O�D
���UI_� HP� '& 8e�w@_T���f� R���Bcg�"KLR�O��T0'����7$BUTTr��R RraLUM��\u���ERV�R�QPa@��S1({ Ơ/GEUR&SF���AM)� LP���E��C�)#�S�1�c�1��P�0�5.�6.�7.�8 ����a@���%j�Q�AS�'R��USR�4) <$Z0� UB�AI΀@�FOC�Q@PRI�Ρm`�� TRI}P�m�UN$ 
5$*	@t�$ kc�j�HR���� q+a��� �G \�0�1���\OS�qAR��V�H�QS1,�?��3�>��� �HU�S1-�����NHOFF!PT0.[p��O' 1,�09-�0GUN?_WIDTH���B_SUB�"p0�'SRT� �/��vA̗` �OR`�RA�U��T����VsCC�М�0 �aC36MFB124� ��/0.D1Gh %bTq���4�.��c)�C�`	%D�RIV���_V�u�,$(��@D��MY_UBY��$V�vA �� B�tC�#�QtBi0hpp+��"L7�BM�1�$��DEY!�E�XG�n��Q_MU���X�10orbҲ�G>ðPACIN΁}�RGC�52�2�32���!RE{����QF����2�02�/TARG�@P1Rc0˦0�R� �03 9d��_�FLA΀r�	�"N�RE�#SW0_A1 �@�!��O���A���3�E���UB�a �\V�HKG�4���:`����05�!CEA���+GWOR!P�5r���MRCV�5 U���OS�M!PC2S�	hB`3hBREF F�FqF\A�0�࿣�0 ��mJ�A~J�A�K�EqFO_RC,KXEKV��S���']#������6 �$���1p؄��b%�pROU�x[2��# 1z5
2�2�P$���� �΀�3��2���Kq�SUL��4;r��6�5� �P@�3�cN�@f��f��c�PL�#�5e�#5e��Ag���|$��70 &�Ôǡ4� ��C�`+�LO�A�d�a� �iu��`�ܓC�pMI��FR��hTj��fR[$HO�h��r�`COMM'#��OB�v{X����؇VP]2�Hq_'SZ3cQu6/cQu12��Nx0Lx�`Lx�WA�eMP�zFA�I�`GT�`AD<�y�!IMRE~T�r_�GP��� ��&ASYNBUF�&VRTD���qσ�OL��D_�:�W:�P�ETU�#�`yQ�0�ECCUP8�VEM:0�e���gV'IRC�q2��le��8u��0CKLAS~^	�VLEX�J�9/������	�LDLDE�F�I<� �r�������Tp�Q��:��
��T1�'������V�� ;``��L���{,�"UR�3�0_R�p󔟑�!� ��U3�/�/�$�`7����0Ғ �TI�Q��SCO�� �Cz�4; #6;�;�;!�;�/�//%*ᢕ���Dx�SЧ@ U_��M<)���JL*��%��q�=)�G�eLIN����W�@XSGAq�> Q ��N�BPK�cH���HOL��  `_�ZABC}?v2�`�XS�@
  ��_ZMPCF}@<�d��?��l!LNI��΀
성� ~A ����q+@��CMC�M0CKsCART�_ٱ#�P_�� $J����������S��S��2UX9W� ��UXE�!A�<��9��d�J�\ɸJ�l���ZPץB� ��b"���Y:!�D" Ca⣖��IGH&3G�?q(!�!��Ap��>�D � T��A�~�$B�PK�'E@K�_a�	c�RV�`F8��Ba�OVCY��@��TU�O0��j�
R�I��1uD��TRA�CEx�V
1^�͐P�HER��E ,�!�������<�$T�b� 2������ �d ��?� �	 HD)uˀ� (�H��0��/d(�$�BTY���O�Z�$�333.x���<�|Z�\�&�8:����C���� CA?��C@�����θ�v2pP��N�2�6���sz����	z���@����� ������&C n��p��	�V3.00�	�rb21�	*�� ����
fffjtW�\p	 ��   ?���Cz�_f�x�� �� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?O��	 O2OO ^OlI0pO�ODlO�O �Kz�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>PbO>O �JO���O��O� (��O0�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯t� ��.��B��v�舿���J�� v��  f+���2f�G����	2 ?�*�c�Nχ�rϫϖ� ���������)��M� 8�q�\�nߧߒ��߶� �������#�I�4�m�@X��|�������� ������8�#�\�G� ��k������������� ��"XC|� ��I�s����� !E3UWi� �������/ A///e/S/�/w/�/�/ �/�/�/?�/+??O? a?k��p?�?�?>?�? �?�?�?�?OOBO0O fOxO�O�OZO�O�O�O �O�O_,_>_�O
_t_ b_�_�_�_�_�_�_�_ oo:o(o^oLo�opo �o�o�o�o�o �o$ H6X~l�� �����?�&��? �h�V���z������� �ԏ
��.����d� R���v�����П⟜� �����*�`�N��� r�����̯��ܯ�� &��J�8�n�\�~��� ��ȿ���ڿ���4� "�D�j�Xώ��:��� ��tϢ�����0��T� B�x�fߜ߮����ߐ� �������P�b�t� ��@���������� ���L�:�p�^��� ������������  6$ZHjl~� ����� 2�� J\n���� ���/
/@/R/d/ v/4/�/�/�/�/�/�/ ??�/<?*?L?r?`? �?�?�?�?�?�?�?�? O8O&O\OJO�OnO�O �O�O�O�O�O�O"__ F_4_V_X_j_�_�_�_ �_p�_ o�_�_Bo0o foTo�oxo�o�o�o�o �o�o,<bP ����v��� �(��8�^�L���p� ����ʏ��ڏ܏�$� �H�6�l�Z���~��� Ɵ���؟���2� � B�h�o������N�ԯ ¯����.��R�@� v�������j�п���� ��*�<�N��^�`� rϨϖ��Ϻ������ �$�J�8�n�\ߒ߀� �ߤ����������4� "�X�F�|�j���� ���������$�6��� V�x�f����������� ����,>��NP�b����  � � �����$TBJOP_�GRP 2W���� ?���C�	�E�� ������X��y�^� �,X�� @� ?����D)̴C2
C랔���wE�{�,d���<-�"z��<p�S�>�g��?#g)? g��B��QBo�'/2'���j/�|%<?D!?���?L�#C  B�Z'�/:/L/^/܀/4H��2/d�;�ŗ-C?��B����/Q?�Cd6����C�p��.v2p��6�?�'�;����CA�?:��?m4��1C�{�CH`R?�?d?�v?�6l4O�6;��?)�2 ?S��PACE�C	���?qO�?O B�E�O�7Kl��2333�?fff?Y-Z�@rO�O�;�%_�' 4__,_Z_�_f_ _�_ �_�_�_�_o�_�_:o@To>oLozo�o~D����!��%	V3.�001rb21�*�`��w� F�� F��. G
� G�(� GG� G�gs G�� G��v G�^ G����G�@�G��; G쑀G��C�H	(�H�� H��H�&��H1�H�;y� r?� F�M4 Fj0 F��` F�v F��V F� G�> G7� G�Zj G�l G����G���G��� G�� G����HS@H���H0) H�B�@=� <��U��l>� V� ^@jQ����
�?�  ��oK�y�� `�\�n���� G����ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �ߪ y���߬߮ !p ���(�:���^�p�� ����	������ j�)�����u�?��� ���������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O���߳O��S��O_ _�O�OK_]_o_�_�_ �_��_����_1�Y� #og�y�ko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i��O�O���O7_ տ�����Ϳ/�A�S� e�wω��_���_�_������$TCPPACTSW  e����I�R e{�#�CH  ��SPEED �2� C�e�  ��5D����_�CFG 	2�D#Ѵ���!Ү��/_SPD��
�>����
�#�:�o®��������NU�Mд���
��OU�T 2��
   ����t��n���� ����������/�"�S��F�X�j�|��ZERO��  ���F�ESTPARS��#����HR��AB_LE 1����R���ٔ�����Q���Ѯ���	���
����������4���RDI��<�&8J\�O����H0��S��� �
 �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?����� z�w���Yk}������n2/� *2�P`�0 3�4�L���2�A@���`�IMEBF_�TT���5��&ќCV�ER2�!ѯF�ќ@R7 1�8ﴰ��d� ��H�7a�6����O�1+�W� DP �[°�,_��O ʱ0[�\_��Y��� 	��^Ĕ_�Y�	�	�P�^��_i W(��P�^�o~������_��$_���\`��`o�to���x7��oɬo�i�5�; 
�o���oEB����\`�L\�<o��������	w!�Q�t��i4�\���wyU͌�0߯� �pL\�DT~�n���L\��N��S_E�V�4��z�T�R�l�~����Ҥ�����Vӌ܏F�T_�������a93�3�E����h�z���� �q�������������u?��"���_[/�Y�k��'��������p*B��ί����������g�9�K���1�`�r�L�w���P���D.�!�@�� �MI_CHAN�G� 
�DBGLVL�G���ETHE�RAD ?���i����0r�:e�u�4:33:9b/:f1 r�2��5�ʆ�4P�RP��@!���!������SNMASK^���o��255.$�0ෳ#�5�G� �OOL?OFS_DI����L�ORQCTRL' �ɦ3�:��5�T��������0� B�T�f�x������ ����������;�*��_���PE_DET�AI<ȉָAPGL�_CONFIG �WIgA�?/�cell/$CID$/grp1c�?�c����������2(]o���4��3���)���40ew ���<����� / /2/�V/h/z/�/ �/�/?/�/�/�/
?? .?�/�/d?v?�?�?�?�?���}S?�?OO8*O<ONO  O�uOTN�R?�O�O�O�O�O _L?)_;_M___q_�_ _�_�_�_�_�_oo �_7oIo[omoo�o o �o�o�o�o�o�o3 EWi{��.� ������A�S� e�w�����*���я� ����+���O�a�s� ������8�͟ߟ�� �'���K�]�o������������Us�er View ���}}1234567890������0�B�J�Ӱ��j���ΩK	�?����Ͽ��� e�w�բ�	�� _�qσϕϧϹ��*� ��SN��%�7�I�[�m����ψ�5�ϼ��߀������u�7�}�6 ��p�������)���}�7_�$�6�H�Z� l�~����}�8��� ���� 2��SY� lCamera٪���� �����BE� .@�Zl~�����  r���/ /(/:/L/^/�/�/ �/��/�/�/ ??$?K�rBɻ/p?�?�? �?�?�?q/�? OO]? 6OHOZOlO~O�O7?I7 ��'O�O�O __$_6_ �?Z_l_~_�O�_�_�_ �_�_�_�OI7��_Jo \ono�o�o�oK_�o�o �o7o"4FXj os^��o���� ���o2�D�V��z� ������ԏ{I7� k� �2�D�V�h�z�!� ��������
�� .�@��I7��ן���� ��¯ԯ母�
��.� y�R�d�v�������S�e�98�����#�5� G��X�}Ϗ�6�����@�������߮�	t0��Z�l�~ߐߢߴ� [������ߣ� �2�D� V�h�z�!�3�y {� ������	��-���Q� c�u������������ ����t���?Qc u��@����, );M_@� S;������/ �)/;/M/�q/�/�/ �/�/�/r��Kb/? )?;?M?_?q?/�?�? �??�?�?OO%O7O �/�+k�?�O�O�O�O �O�O�?__%_pOI_ [_m__�_�_JO��{ :_�_oo%o7oIo�O moo�o�_�o�o�o�ox�o�]  �Y >Pbt���������    :�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d��v��  
�`( � �2p( 	 �������ο�� (��8�:�Lς�pϦ����ϐ�$� � ^o�!�3ߦoW�i�{� �ߟ߱߸S�������� F�#�5�G�Y�k�}��� ������������ 1�C���g�y������ ��������	P�b�? Qc������� �()pM_ q������� 6/%/7/I/[/m/� ��/�/�//�/�/? !?3?E?�/i?{?�?�/ �?�?�?�?�?OR?/O AOSO�?wO�O�O�O�O �OO*O__+_rOO_ a_s_�_�_�_�O�_�_ �_8_o'o9oKo]ooo �_�o�o�o�_�o�o�o #5|o�ok}� �o������T 1�C�U��y������� ��ӏ���	��b�?��Q�c�u���������@� ��ȟڟ쟻������)frh�:\tpgl\r�obots\r2�000ix&�b_�210f.xml ��P�b�t����������ί���� �dummy"�;�?�Q� c�u���������Ͽ� �
��.�;�M�_�q� �ϕϧϹ�������� �*�7�I�[�m�ߑ�@�ߵ����������� �)�;�M�_�q��� ������������%� 7�I�[�m�������� ��������!3E Wi{����� ���/ASe w��������;� �8?8�?��"/ �/@/B/T/v/�/�/ �/�/�/�/?�/?B?�,?N?x?b?�?�?�;��$TPGL_OUTPUT �   ?O���3;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__Б_�_�3 �@23�45678901 �_�_�_�_o o(c� �_Ooaoso�o�o�oAo��o�o�o'�j} 1Yk}��9K �����1��?� g�y�������G���� ��	��-�ŏ׏c�u� ��������U�˟�� �)�;�ӟI�q����� ����Q�c����%� 7�I��W�������� ǿ_�տ���!�3�E� ݿ�{ύϟϱ����� m�����/�A�S��� a߉ߛ߭߿���i�A}!��+�=�O�a��r�@/���* ( 	 �_���� ���%��I�7�Y�[� m������������� ��E3iW�{ ������/�V� "7ewS ������RP
/ /�@/R/0/v/�/� �/�/`/�/�/�/�/*? <?�/`?r??�?�?�? �?�?H?�?O�?OJO \O:O�O�O�?�O�OjO �O�O�O"_4_�O _j_ |__�_�_�_�_�_R_ oo�_BoTo2odo�o �_o�o�oto�o�o ,>�obt�� ���J\�(�� L�^�<��������ʏ l�ڏ �ޏ��6�H��� l�~� �������؟� T��� ��V�h�F� �����¯ԯv���
� �.�@���,�v���*��������������$�TPOFF_LI�M K|�ӱ��|��N_S]V�  x�%�� �P_MON CG�*�|��2x��STRTC�HK CE���M�VTCOMP�AT:���I�VWV_AR Z��Ȗh��� ��|��m��_DEFP�ROG %��%�FOLGE01�1ߢ�_DISP�LAY���/�IN�ST_MSK  �� k�INU�SER��-�LCK��܊�QUICKM�EN��q�SCRE��C��t_scq���!�&�%��7�ST��E�RAC�E_CFG �Z����	�
�?���HNL 2E��#���� � �������"�4�F�X��j���ITEM 2��� �%$1�23456789y0����  =<��x������  !�����Jӫ�k �����); _�/U��� �	�7�	// ?/���A/��/ �/�/3/�/W/i/{/�/ M?�/q?�?�/�??? �?A?Oe?%O7O�?MO �?O�O�?�OO�O�O �OaO	_�O�O�O#_�O y_�_�__�_9_K_]_ �_�_�_Soeo�_qo�_ �_�o#o�oGo}o /�o�o|�o��o� �SCUg��� �[���������-� ?���c��5�G���S� Ϗ��w�ş)���� _������^���y�ݟ �����ů7����m� -���=�c�u�ٯ���� �!���E���)ύ� Mϱ�ÿտY�q���� ��A���e�w�@ߛ�[� ��ߑ��ϧ��+���ʀ�S����F��g  u�F� ��P�F�
 ]��j����(�UD1:\������R_GR�P 1 ��� 	 @P�������1��U�C�y�g�� �����s����������?�  ) I7m[��� ����3!WEg�	�ա� q��m�/�'//7/ ]/���/���/���/ �k�/#??G?5?k? Y?�?}?�?�?�?�?�? O�?1OOAO���O ��Oe/�O�O�O	_�O -_k/Q_�/x_�/u_�_ QO�_MO�_�_oo'o Mo;oqo_o�o�o�o�o �o�o�o7uOS e#_�_���� ��M_3��_Z��_~� �_����ՏÏ��� ��A�/�Q�S�e��� �������џ�Eo�5�G��SCB 2!� ������ ����ϯ�������X_SCREEN� 1"��
 �}�ipnl/X�g?en.htm$�w����������P�P�anel set�upü}	ind?ex.STMÿ���1�C�U�̷
Ro�bot Info e�9�ϱ��������� �τ�1�C� U�g�yߋ�߯�&��� ����	��-�߶�c� u�����4�b�X� ��)�;�M�_���� �����������x� ��7I[m� 6,���!3��W3�UALRM_MSG ?D��Q� RD�� ����/
//:/�@/q/d/�/�/�/mS�EV  {��&kECFG �$e�  D7�A�1   B�N+N�Q�0�4� � A aX��2?F0�4=�XxF0jb?_KX��lz?a�X�[��?^�0S�?k_h�0v�?^��0���?�0��?_�X���!GR�P 2%e� 0�*0�2�p������5r?��>Vvտ�FN/?͇��,��&0 v��On��O�O�O�Oj�I_DEFPRO�w+F� (%�MAKRO050� .(_-Q00343  _/_05CP�/ _Nm_�_�_�_�_�_��_o�_#oHo�DINUSER  ]��ONoI_MENH�IST 1&e� � ( P���-/SOFTP�ART/GENL�INK?curr�ent=edit�page,FOLGE125,1�o�&D�o�o�c011,jPv����;y%HZ~�`np20 s��,�7}'�Zuomenu�b37�o ��������C�gw�p v��#�5�Č+ԏ��UP024,20�D�������?�Y�c�98���$�6�H�ן��a71��a�������Ы�6a�a6o���  �2�D�V�̓므��� ����ȿڿi����"� 4�F�X��|ώϠϲ� ����e�w���0�B� T�f��ϊߜ߮����� ��s���,�>�P�b� ������������ ݯ�(�:�L�^�p��� ����������� �� $6HZl~� ������2 DVhz��� ���
/�./@/R/ d/v/�/�/)/�/�/�/ �/??�<?N?`?r? �?�?�?�/�?�?�?O O&O�?JO\OnO�O�O �O3O�O�O�O�O_"_ 4_�OX_j_|_�_�_�_ A_�_�_�_oo0o�_ Tofoxo�o�o�o�oOo �o�o,>)?�o t������o� ��(�:�L��p��� ������ʏY�k� �� $�6�H�Z��~����� ��Ɵ؟g���� �2� D�V����������¯ ԯ�u�
��.�@�R��d�Oz�$UI_P�ANEDATA �1(������  	��}/frh/c�gtp/wide�dev.stm �&C1=OFF&�B2=Save&�ACTION=101&C2=8p������ )prsim�<�  }?��c�uχϙϫϽ� ) ���������+�=�$� a�H߅ߗ�~߻ߢ���p�����Lv�[q�7�JǨ�vagmn1��*�m������ual����O� � �$�6�H�Z��~�e� �������������� 2V=z�s�#� �������� ,>P�t�� �����Y/(/ /L/3/p/�/i/�/�/ �/�/�/ ?�/$??H? Z?���?�?�?�?�? �?=?O�2ODOVOhO zO�O�OO�O�O�O�O 
___@_'_d_v_]_ �_�_�_�_�_�_g?y? *o<oNo`oro�o�_�o �o-O�o�o&8 �o\C��y�� �����4�F�-� j�Q���oo�o֏� ����0���T��ox� ��������ҟ9���� �,��P�b�I���m� ����ί�ǯ��(� :�����p��������� ʿ��a��$�6�H� Z�l�~�忢ω��ϭ� ������ ��D�V�=� z�aߞ߰ߗ���G�Y� 
��.�@�R�d�߈� ��Ͼ��������� �<�#�`�r�Y���}� ����������&`J1n����}�@���� )� 7��&cu��� �$��/��;/ "/_/F/�/�/|/�/�/��/�/�/?��������$UI_POST�YPE  ���� 	 ��?��E2QUI�CKMEN  �T;c7�?�8RESTORE 1)���  �?���?�3�?��mODOVOhOzO�O /O�O�O�O�O�O�O_ ._@_R_d_Oq_�_�_ _�_�_�_oo�_<o No`oro�o�o9o�o�o �o�o�_!3�o n����Y�� ��"��F�X�j�|� ��9C�����1��� �0�B�T���x����� ����c������,� ׏9�K�]�ϟ������ ί௃���(�:�L� ^����������ʿ�7oSCRE�0?�=u1sc�0Wu2�3�4�U5�6�7�8�E2USER����Sks�f�3f�4f�U5f�6f�7f�8f��E0NDO_CFG� *T;� �E0P�DATE P���KS_24��1G�_INFO �1+�����10%�FOLGE01�1п�� ��% �Eߣ�3�t�Wߘߪ� �����������(�:���^�p���OFFS_ET .�=q� l��0s���������� �!�N�E�W���[��� ����������/y��?{
c2����t�SEUFRAM/E  d������RTOL_ABRqT����ENB�~�GRP 1/�9��1Cz  A� :8l�8J\n�B����
�0U����MSK  h���	N�%���%KH/�2VCCMf��0��]"MR {26T9 d��¼�	��m2%~?XC56 *�/�&�X���0�5���A@�p��L.-�k7?d�7?I?�v?�!q?�?5�A��l��?�?l�� B����1l��5�?O b??OOcONO�OrO�O �O�O�O8O�O___ M_ Oq_�_d��!�!�/ �_�/�/�/??'?o �O\oSo1_�o�o�?�? �o�?__�o"io{o= jU�y���- ���	�B�U_f�x� ����!�_���_�_�_ oo'o��\�S�1� �����o�oڟ�o_��� "�i�{�=�j�U���y� ����֯-���ɯ�	� B�U�f�x����=��� ��͏ߏ���'�� �\�S�1��ϤϷ�ɟ ���_���"�i�{�=� j�Uߎ�y߲ߝ���-� �����	�B�U�f�x��O/ISIONTM�OU� $r%����d#7�K ��LT/ F�R:\��\DAT�A\�� �� wMC��LOG��   UD1���EX��' ?B@ ��O� ��7/m� �q���� ��  =	 �1- n6  G-��T�L�&,��<���=�����T����TRAIAN6������"8�+ (:���S.�S as��������'9KX&L�EXE��9�+�!1�-eR,MPHASOE  k%�#�R�]!SHIFTME�NU 1:�+
 �<\�6//���� �!/Z/1/C/�/g/y/ �/�/�/�/?�/�/D?�?-?z?Q?	LIVE/SNAPn3vsfliv���?^3�� SETyU�0�2menu�?��?d?)O;OB��;����	(H'O�Oh\����� ��@⹭A�B8`�`��������A�B��C���G ��KSFME��0����� �M�O�<��z��W�AITDINEN�D���Q@WOK C �X[]��w_S�_�^YTIM�����\GH_�]j_�[�_�Z�_�Z�_\XRELE��gU@T����AS_ACT�0
h�aq����d�� =���b%$FOLGE�011.	r00�0���dRDIS��0�oAPV_AXSMRG`2>bJ<��O���Gp4 _IR  ��᥀����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z�����oZABC31?bI&�� ,�=�2��ܬ ¯�����
��Y����MPCF_G 1@S}0A�������ҿ�������,�b�MPz��AbI  �@���:��Q8�|O����t��Ϙ�?� T�������D����k�-ߞ߰��ѿp����� ������	�l�E��i� {�ߟ�R�\�n߀ߚ� �����2���e�w�� ��������.�� d�=OZ�s�@�� \�����'9 ����Tf���� �&�/5/� \//�/B/T/f/x/�/ �/F��(?:?L?v>ȣ�u�(PBS{j�P_�CYLINDERw 2CS{ ��& ,(  *�?��=�#�?O�?8OM �/nO�O�N�?�O$O �O�O�O_RO3_E_W_ �O{__�O�_�_�_�_`*_oof�R�2DSw�`�P�"�hoxl�s�/��o�o�o��o�o�1�qA��o*yo�o` �o��o}�	�� ?y&�uJ��Z��� �m����?��׏��_�4�F����2SPH�ERE 2E�=� o_���_��͟����_ L�'�9�i_]���⟓� z���������F�X� 5���Y�@�R���֯���ſ׿N�ZZ  �$��4