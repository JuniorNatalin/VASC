��   2W�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���C�ELL_GRP_�T   � �$'FRAME �$MOUN�T_LOCCCF�_METHOD � $CPY_SRC_IDX_�PLATFRM_�OFSCtDIM~_ $BASE{ �FSETC��A�UX_ORDER�   �X�YZ_MAP �� �LEN�GTH�TTCH�_GP_M~ a AUTORAIL_���$$CLA�SS  ��i���D��D�8LOOR ���D8�?���O��/, � 1 F �H8=_`_��D'�82 �����K!/3/E//i/{/�-_ �/�/�/pO,��p 8!�/ �/?/g?y?�?]?�? �?�?�/�?�?�?�/C?E?�13OEOWOY?�O �O�O�O�O	__	O3_@E__1O�O�O�A{_ �_�_�O�_	oo�_?o�QocoQ_{o�ogo�$�MNU>A�R�d  8K�_�_ ��o	=?Q s������	� ��?�)�K�u�_��� �������ˏݏ�� �5�7�I�k������ ˟��ן���7�!� C�m�W�y�������ٯ ïկ����b!�K� 2�G�i�k�}���ɿ�� տ����5��A�k� U�wϡϋϭ������� ���	�C�-�?�a�c� uߗ��߫�������� -��9�c�M�o��� �����������;� %�7�Y�[�A�1q��� ����������- 9cMo���� ���;%G q[m����� ��%//1/[/E/g/ �/{/�/�/�/�/�/�/ 	?3????i?S?e?�? �?�?�?�?��A�?O �?O1O3OEOgO�O{O �O�O�O�O�O�O	_3_ _?_i_S_u_�_�_�_ �_�_�_o�_o)o+o =o_o�oso�o�o�o�o �o�o+7aK m����������!�#�  �$�MNUFRAME�NUM  W�>�X�D � k�TOOL ?A��������\ @��;�.L�K��L������3��Ł'	��D�;s3��C�zff��5��?�W���O��j�� C���C L��Y�[�#�E�o�Y� {�������۟ş�� ���G�1�S�}�g��� �������ӯ��	� �=�g�Q�s������� ӿ��߿	���?�)� K�u�_ρϫϕϧ��� ��������5�_�I� kߕ�ߡ��ߵ���� ���7�!�C�m�W�y� �������ﱂp��� ��n�2�4�F�h���|� ������������
4 @jTv��� �����*, >`�t���� ��/,//8/b/L/ n/�/�/�/�/�/�/�/ �/ ?"?$?6?X?�?l? �?�?�?�?�?�?�?$O O0OZODOfO�OzO�O �O�O�O�O�O�O__
�13_q_X_m_�_�_ �_�_�_�_�_%oo1o [oEogo�o{o�o�o�o �o�o�o	3/i Se������ ���)�S�=�_��� s�������ˏ��ߏ� +��'�a�K�]���� ����ߟɟ����!� K�5�W���k������� ï�ׯ��#���Y� C�U�w�y��A��Ϳ ��ɿ����!�K�5� Wρ�kύϷϡ����� ����#��/�Y�C�e� ��yߋ��߯������� ���C�-�O�y�c�� ������������ '�Q�;�]���q����� ����������;% Gq[}���� ���I3U i{������  �$MNUT�OOLNUM  �
 
 ?D  @!