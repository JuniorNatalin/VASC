��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �
  ����
��WVAMP_T �  $X�1  $X2�AY@h/FC~5  $2�ENBA $DTo  / _R2� d ENAB�LEDnSCHD�_NUMA  ��/ CFG5�� $GROUP��$z ACCEL�@�G$MAX�_FREQ�2 L��DWEL�DE�BUG�PREW�SOUT�P�ULSEASHsIFt 7TYP4�$USE_AE�F} 4$GDO��  f0 �r?�NpWE�AVE_TSK u�V�_GP��SUPPORT_�CFnCNVT_?DONE p }�k}GRP 2�r�� _� �}$� TIME1�to$2'EXT� �(1#&(MODE_�SW�CO3 SW�IT � X/ PH�AX6  4 �� ECC$�T�ERMNnPE�AKno!AL � \ � �!I֑$�!N_VSTAR�#!r"ؾ�"�%�CY�CL42 ��/ � Tv"b $�CUR_REL_܂ �! x/ WP�R5 � 
$wCEN� _RI3_RADIU��XIz ] ZI�MUTi!$ELEVATIONg5�� N�CONTI�NUOe2q �ME�XAC=PE�qt1�6  H~ >�UENCYA��ITUD4�2RI�GHC�2LEBL�_ANG1 ��OTF_� 	�  $3A�b�ET��n3C!�$ORGjHFSBKjH��P��C\��DLDW�HR�E�_�3�B�C��D�B��C�@�D�A�CCHG��G	Q�F	Q�F	Q�FINC�G=Q�F=Q�F=Q��F�AVCPYC� _�T�\#�Y~P#�@S�Y��H)@�UP�D"0n�$$C�LASS  �����Q��8 �P��� VA2�U�� �   =?��@�  aa �U�To-o?oQoco�P��TN 2 �[ �f��ue@O�i�oc�Q� � F�Ua	`��`�d\ �` �����=������b ����.pqUcw -�ut(q��uvp�P���xu��d�aPq��&�8���0�q,B��}a� u s�s�a� s�������֏b�Q� w 2�[
Ta�SI��}�v���F� ,�?1�'��P�0��P�P�a ��0�l�jk��ҟ������,�>�ll�FIGURE 8��3�:�a0�*�X� e�ۯү�������L�R�d�v������T�CIR1q� dֿA���B�,�>���0�����:�`�B���ϲ�������nj� pq�(qG�V�E�@�����`+ݳ� �ߗߩ߻����������'�9�S�Lp��%��B�5)�� T�`���p���䏟 ��w��#�5�G�Y�k��}���mkTr?ianglej��� >�,߂�L���D�Q cu������� �������X� +X2D���� �//'/9/�} ,>l/�/���/ ?!?3?E?W?i?{?�?��C��?nhE��? �?OO,O>OPObOtO �O�O�O�O�O�O�K�? �O�?�?H_Z_l_~_�_ �_�_�_�_�_�_o o�2o|mSCHEXT?ENB  ��c��STATE 2�k @o�o�o��o�oNgWPR ����}��_O�TF 	�oa�@ � qq]qQcuv�qu�A�os�u@�  <#�
�?��^��1u_GP 2;| �Io(�:��� �����e+