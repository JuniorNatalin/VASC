A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �PNIO_AN_T   L $AO_ADR  $AO_SHIFT  $AO_VALID  $AI_ADR  $AI_SHIFT  $AI_VALID   �PNIO_CFG_T � �$VERSION $COMMENT $CUSTOM  $CUSTOM2  $DEV_ENB  $CON_ENB  $TMP  $START_MODE  $NUM_LST  $NUM_MOD  $CHG_DIG_PRT  $PS_MAX_DIG_   $MAX_DIG_PRT  $C_DI_PRT  $C_DO_PRT  $C_AI_PRT  $C_AO_PRT  $C_WI_PRT  $C_WO_PRT  $C_WSTI_PRT  $C_WSTO_PRT  $C_DI_OFS  $C_DO_OFS  $C_AI_OFS  $C_AO_OFS  $C_WI_OFS  $C_WO_OFS  $C_WSTI_OFS  $C_WSTO_OFS  $D_DI_PRT  $D_DO_PRT  $D_AI_PRT  $D_AO_PRT  $C_HOLD_DI  $D_HOLD_DI  $ACT_INDEX  $ACT_OPCODE  $ACK_INDEX  $ACK_OPCODE  $INIT_PRM  $ANNOT_NAME $ANNOT_ORDER $ANNOT_HW  $ANNOT_REV  $ANNOT_SW1  $ANNOT_SW2  $ANNOT_SW3  $DEV_SLOT  $DEV_VID  $DEV_DID  $DEV_INST  $PS_CP16XX_W   $CP16XX_W1  $CP16XX_W2  $CP16XX_W3  $CP16XX_PK1  $CP16XX_PK2  $DEV_SEARCH  $DEV_COMCHK  $TP_WAIT_ACT  $PG_WAIT_ACT  $MAIN_REQ  $MAIN_PARAM  $MAIN_EXEC  $CON_ER1SHOT  $DEV_ER1SHOT  $ENABLE_WIO  $ASG_UOP  $WD_TIME  $WD_ENABLE  $TP_DEBUG  $SCAN_TIME  $D_DEFAULT  $PG_WAIT_ST  $DEV_APDU  $PWRCLR1SHOT  $COMCLR1SHOT  $CON_IOCLR1  $CON_IOCLR2  $DEV_IOCLR1  $DEV_IOCLR2  $FLAG  $AUTO_OPMODE  $PWOFF_ALARM  $ERRDEACT_I  $ENB_DEVCHK1  $ENB_DEVCHK2  $INIT_DEVCHK  $CYC_DEVCHK  $CYC_IOSTAT  $BOARD_SV  $WD_SV  $DEV_OP_SV  $DEV_ABO_SV  $DEV_OFF_SV  $DEV_MIS_SV  $CON_OP_SV  $CON_ALM_SV  $CON_OFF_SV  $CON_CLR_SV  $TIMEO_SV  $DEV_MOD_SV  $DEV_SMD_SV  $CON_CFG_SV  $DEV_DACT_SV  $DEV_STOP_SV  $CON_STOP_SV  $CON_NOPR_SV  $READIN_SV  $PWOFF_SV  $AUTO_OP_SV  $ALARM1_SV  $ALARM2_SV  $ALARM3_SV  $UPDATE  $TRC_FILE $TRC_MAXSIZE  $TRC_ENABLE  $TRC_TIME  $TRC_DEST  $TRC_DEPTH  $TRC_GROUP  $TRC_OUT  $ULONG1  $ULONG2  $ULONG3  $ULONG4  $ULONG5  $ULONG6  $ULONG7  $ULONG8  $UBYTE1  $UBYTE2  $UBYTE3  $UBYTE4  $UBYTE5  $UBYTE6  $UBYTE7  $UBYTE8  $UBYTE9  $UBYTE10  $UBYTE11  $UBYTE12  $UBYTE13  $UBYTE14  $UBYTE15  $UBYTE16  $UBYTE17  $UBYTE18  $UBYTE19  $UBYTE20  ,�PNIO_CFG2_T  ($VER_INFO $COMMENT $DIV_DELTA  $DIV_ENB  $CON_OPTION  $DEV_OPTION  $IOR_TRANS  $IOR_OPTION  $RST_CONT  $RST_RESET  $RST_CYCLIC  $RST_SEV  $RST_INTVL  $PS_PS_MOD_L   $PS_MOD_LOW  $PS_MOD_HI  $OPT1_SEV  $OPT2_SEV  $USHORT1  $USHORT2  $USHORT3  $USHORT4  $USHORT5  $USHORT6  $USHORT7  $USHORT8  $USHORT9  $USHORT10  $USHORT11  $USHORT12  $USHORT13  $USHORT14  $USHORT15  $USHORT16  $USHORT17  $USHORT18  $USHORT19  $FW_VER_REQ   $FW_VER_STOP  $UNCFIRM_SEV   4�PNIO_DB_T  � $COMMENT $BASE_MODID  $IO_MOD1  $I_MOD1  $O_MOD1  $IO_MOD4  $I_MOD4  $O_MOD4  $IO_MOD16  $I_MOD16  $O_MOD16  $IO_MOD20  $I_MOD20  $O_MOD20  $IO_MOD64  $I_MOD64  $O_MOD64  $ULONG1  $ULONG2  $ULONG3  �PNIO_DBG_T  � $START_REPWR  $START_TIMED  $DELAY_TIME  $ULONG1  $ULONG2  $ULONG3  $ULONG4  $ULONG5  $ULONG6  $ULONG7  $ULONG8  $ADDR1  $ADDR2  $ADDR3  $ADDR4  $ADDR5  $ADDR6  $ADDR7  $ADDR8  �PNIO_DIAG_T  � $FW_VERSION !$CNTR_STAT  $DEV_STAT  $DRIVER_STAT  $PROC1_STAT  $PROC2_STAT  $PROC3_STAT  $CON_I_STAT  $CON_O_STAT  $ULONG1  $ULONG2  $ULONG3  $ULONG4  $ULONG5  $ULONG6  $ULONG7  $ULONG8  L�PNIO_DIAG2_T  A$ST_NAME1 �$ST_NAME2 �$ST_TYPE1 �$ST_TYPE2 �$IP_ADDR !$IP_MASK !$ROUTER !$ALM_MSG1 =$ALM_MSG2 =$ALM_POST  $ALM_SEV  $ALM_OPTION  $STORM_RESET  $STORM_ST  $STORM_UNKST  $STORM_EXIST  $CMD_BUSY  $CMD_TYPE  $CMD_REQ  $CMD_ACK  $CMD_INFO  $BACKUP_STAT  $CONFIG_STAT  $FWV !$SNR !$HWV  $R1  $R2  $CP_STATE  $EXT_PAR  $MAC !$MLFB !$F_IP !$F_MASK !$F_GW_IP !$PS_R3_1   $R3_1  $R3_2  $SDB_COUNT  $DAP_SLOT  $MODID   $TIME1  $TIME2  $TIME3  $TIME4  $TIME5  $TIME6  $TIME7  $TIME8  $MONITOR1  $MONITOR2  $MONITOR3  $MONITOR4  $MONITOR5  $MONITOR6  $MONITOR7  $MONITOR8  $STATUS1  $STATUS2  $STATUS3  $STATUS4  $STATUS5  $STATUS6  $STATUS7  $STATUS8  �PNIO_DL_T  � $PATH_XDB A$PATH_FIRM A$TIMEO_XDB  $TIMEO_FIRM  $OPCODE_XDB  $OPCODE_FIRM  $NO_FIRM_ST  $XDB_SEV  $FIRM_SEV  $DOWNLOAD  $WAIT_RATIO1  $WAIT_RATIO2   \�PNIO_DL2_T l u$ST_TYPE1 �$ST_TYPE2 �$BACK_XDB A$BACK_FIRM A$BACK_SNUM A$K_BACKUP  $K_DOWNLOAD  $K_OPERATION  $FLAG_BACKUP  $FLAG_CHECK  $COLD_FLAG  $COLD_TIMEO  $COLD_TIME2  $TIMEO_BXDB  $TIME2_BXDB  $CPY_BXDB  $BLOCK_BXDB  $WAIT1_BXDB  $WAIT2_BXDB  $SEG_BXDB  $CONF_BXDB  $PRM_BXDB  $PNIO_BXDB1  $PNIO_BXDB2  $PNIO_BXDB3  $PNIO_BXDB4  $TIMEO_BFIRM  $TIME2_BFIRM  $PS_BUFF_BFI   $BUFF_BFIRM  $BLOCK_BFIRM  $WAIT_BFIRM  $CONF_BFIRM  $PRM_BFIRM  $PNIO_BFIRM1  $PNIO_BFIRM2  $PNIO_BFIRM3  $PNIO_BFIRM4  $FILE_BTO  $FILE_DTO1  $FILE_DTO2  $FILE_BSIZE  $FILE_DSIZE  $BXDB_SEV1  $BXDB_SEV2  $BXDB_SEV3  $BXDB_SEV4  $BFIRM_SEV1  $BFIRM_SEV2  $BFIRM_SEV3  $BFIRM_SEV4  $BACKUP_SEV  $XDBMIS_SEV  $XDBCHK_SEV  $BADMOD_SEV  $WNGGSD_SEV  $SETTING_SEV  $SAFE1_SEV  $DOWN_FW_SEV  $OLDBACK_SEV  $DID_SET_SEV  $ALM1_SEV  $ALM2_SEV  $SERVLIB  $LOCK  $PNIO_HI  $PNCM_HI  $PNSV_HI  $PNSV_LO  $PNSV_TIMEO1  $PNSV_TIMEO2  $PNSV_CONFIG  $PNIO_IOC  $PNIO_IOD  $PNIO_START1  $PNIO_START2  $CHECK_BACK  $REMOTE  $HOLD_CMT  $CHECK_FWV  $PS_STORM_EN   $STORM_ENB  $STORM_TIME  $STORM_COUNT  $STORMALM_SV  $STORMCLR_SV  $CYC_ALM  $INIT_PRM1  $INIT_PRM2  $INIT_PRM3  $INIT_PRM4  $INIT_PRM5  $INIT_PRM6  $SYNC_NUM1  $SYNC_NUM2  $SYNC_PRM1  $SYNC_PRM2  $SYNC_PRM3  $SYNC_PRM4  $SYNC_PRM5  $SYNC_PRM6  $OUT_FILE1 $OUT_FILE2 $FLAG1  $FLAG2  $FLAG3  $FLAG4  $FLAG5  $FLAG6  $FLAG7  $FLAG8  $FLAG9  $FLAG10  $FLAG11  $FLAG12  $CLASSCODE1   $CLASSCODE2   �PNIO_LST_T 	 � $COMMENT $ENABLE  $ADDRESS  $LENGTH  $STATION  $SLOT  $SUBSLOT  $ADDRTYPE  $IODATATYPE  $DATATYPE  $COMTYPE  $ERRDEACT  $IN_INDEX  $OUT_INDEX  $CONFIG  $STATUS1  $STATUS2  $STATUS3  �PNIO_IM0_T 
 � $VERH  $VERL  $RES1  $RES2  $VID  $HWR  $SRP  $FE  $BF  $IC  $ORDER_NO $SERIAL_NO $RC  $PI  $PST  $VMA  $VMI  $IMS  $RES3  $RES4   ��PNIO_MOD_T  � 
$COMMENT $SLOT  $SUBSLOT  $MODID  $SUBSLOTID  $NUM_INPUT  $NUM_OUTPUT  $IO_TYPE  $DATA_SIZE  $DATA_TYPE  ��PNIO_WRK_T H $OUT_FILE $OUT_MODE  $DEV_ENB0  $CON_ENB0  $TP_DEBUG  $START_MODE0  $PWOFF_FLAG  $WIO_ENABLE  $CON_FLAG1  $CON_FLAG2  $DEV_FLAG1  $DEV_FLAG2  $COM_FLAG1  $COM_FLAG2  $UBYTE1  $UBYTE2  $PS_PNIO_SYS   $PNIO_SYSV  $ADDR1  $ADDR2  $ADDR3  $ADDR4  $ADDR5  $ADDR6  $ADDR7  $ADDR8  �$$CLASS  ������   N    N�$PNIO_AN 2 ������N�                                                                                                
         
                                                                                                                                                                                                                 "         "         $         $         &         &         (         (         *         *         ,         ,         .         .         0         0       �$PNIO_CFG ������N�V820P02 131028            �                                      �                  @   @  �  �                                  FANUC Robot Controller        A05B-2600-J930              V    �  �     �   d  �  �  �  ���                 �          �,                   mc:pniotrc.txt                                                                                  ��$PNIO_CFG2 ������N��                          �                           @        �                                            �$PNIO_DB 2������N�  hCP1604 DAP V2.6                     !   "   #   $   %   &   '   (   5   6   7   )   0   1     !  "CP1604 DAP V2.6(M)                  !   "   #   $   %   &   '   (   5   6   7   )   0   1     !  "CP1616 DAP V2.6                     !   "   #   $   %   &   '   (   5   6   7   )   0   1     !  "CP1616 DAP V2.6(M)                  !   "   #   $   %   &   '   (   5   6   7   )   0   1     !  "
CP16XX DAP                  ��       !   "   #   $   %   &   '   (   5   6   7   )   0   1     !  "                                                                                                                                                                                                                                                                                                                     �$PNIO_DBG ������N�      �                                                                �$PNIO_DIAG ������N�!2.6.1.0                             �  �                ۑ�ۓ�                                �$PNIO_DIAG2 ������N �kjltvr111120r01rs--kux                                                                                                                �                                                                                                                                       �S7-PC                                                                                                                                 �                                                                                                                                       !172.26.30.220                     !255.255.255.0                     !172.26.30.1                       =                                                               =                                                                                                                     !                                   !                                         !                                   !                                   !                                   !                                   !                                   �                         7   6                                                                                                                                                    �$PNIO_DL ������N�AMC:PCST_1.XDB                                                     AMC:\pn2610.FWL .3.9.FWL l                                          �X         d d�$PNIO_DL2 ������N��FANUC Robot Controller                                                                                                                �                                                                                                                                       AFR:S7PRJ.XDB                                                      AMC:\fw_image.fwl                                                  A�                                                                                         ,X,X            n �  ���  �   �     n �     x��             EEE���            �     ( �   � � � � �                MC:\                      MC:\                                                  �$PNIO_DLST 2	������N   D                                ?�       �                                                       v      �                                                      v      �                                                    ?�       �                                                      ?�       �                                                     �      �                                                     �      �                                                     ?�       �                                                      �      �                                                    �      �                                                     �      �                                                    ?�       �                                                       X   
   �                                                      X   
   �                                                    ?�       �                                                       l   
   �                                                      l   
   �                                                    ?�       �                                                       b      �                                                      b      �                                                    ?�       �                                                      ?�       �                                                      �      �                                                    �      �                                                     �      �                                                    ?�       �                                                       H      �                                                     H      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �$PNIO_IM0 
������N�   � VA05B-2600-J930        F174555                   �$PNIO_LST 2	������N�  D                                ?�       �                                                       v      �                                                      v      �                                                    ?�       �                                                      ?�       �                                                     �      �                                                     �      �                                                     ?�       �                                                      �      �                                                    �      �                                                     �      �                                                    ?�       �                                                       X   
   �                                                      X   
   �                                                    ?�       �                                                       l   
   �                                                      l   
   �                                                    ?�       �                                                       b      �                                                      b      �                                                    ?�       �                                                      ?�       �                                                      �      �                                                    �      �                                                     �      �                                                    ?�       �                                                       H      �                                                     H      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �$PNIO_MOD 2������N�  @DAP V2.6                                                 SAFE 8 BYTE                                              32 BYTE                            7                     32 BYTE                            6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �$PNIO_STM  ������N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �$PNIO_WRK ������N �                                         ����                                