A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DCSS_CPC_T   � $COMMENT $ENABLE  $MODE  $GRP_NUM  $MODEL_NUM   $UFRM_NUM  $NUM_VTX  $X   $Y   $Z1  $Z2  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD  �DCSS_CSC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $TCP  $UFRM_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  �DCSS_GRP_T  � $TCPCHG_SIZE  $APSPD_MODE  $ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $APSPD_JMODE   	$ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$TCP_SEL  H�DCSS_GSTAT_T  D $FP_BASE $LINK_BASE ! 	$LINK_BASE_V ! 	$LINK_BASE_H ! 	 ��DCSS_JPC_T  � $COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $UPR_LIM  $LWR_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $ENBL_CALMD   X�DCSS_JSC_T  | 
$COMMENT $ENABLE  $MODE  $GRP_NUM  $AXS_NUM  $SPD_LIM  $STOP_TYP  $DSBIO_TYP  $DSBIO_IDX  $STOP_TOL  P�DCSS_ELEM_T  T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    p�DCSS_MODEL_T   $COMMENT $ELEM 2 
�DCSS_PSTAT_T  � 	$STATUS_CPC    $STATUS_CSC   $STATUS_JPC   ($STATUS_JSC   ($USER_MODEL   $ROBOT_MODEL   $USER_ELEM   $ROBOT_ELEM   $CUR_TCP   ��DCSS_SETUP_T 	 l $DISP_MGN  $INP_ASSIST  $TOOLCHG_ENB  $DO_TYP  $DO_IDX  $DO_MGN  $CALMD_ENB  $CALMD_STAT  t�DCSS_T1SC_T 
  $ENABLE  $SPD_LIM  �DCSS_TCP_T  l $COMMENT $UTOOL_NUM  $MODEL_NUM  $VRFYIO_TYP  $VRFYIO_IDX  $X  $Y  $Z  $W  $P  $R  ��DCSS_SPH_T  ( $SIZE  $DATA1  $DATA2  $DATA3  �DCSS_BOX_T  8 $SIZE1  $SIZE2  $SIZE3  $X  $Y  $Z  $R  0�DCSS_TUIRO_T  , $TYPE  $SPHERE 2 $BOX $BOX_S 2 @�DCSS_TUIZN_T  0 $ENABLE  $X   $Y   $Z_UPR  $Z_LWR  �DCSS_UFRM_T  @ $COMMENT $UFRM_NUM  $X  $Y  $Z  $W  $P  $R  �$$CLASS  ������   Q    Q�$DCSS_CPC 2 ������Q   ��                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �                                       ����                                                                                                           �$DCSS_CSC 2������Q  D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_GRP 2������Q  �                         	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                                                  	                                      	                                      	                                      	                                      	                                         �$DCSS_GSTAT 2������Q  ,8���n��M|?}�5?�<���=�q��U?~��=���D�+MC�e�D��0��� 	 88�?|b>1�]    �j�4���?�  >1�]�|b4��ZC�0�B��    ���8������?Q���N�8�����>1�]�|b4��Z�d���!Z�DW����8��N������&?�=����Q�z>1�]�|b4��ZB&�p@�>��em���8�>1ώ�|k6�4��N������&?�+=����Q�zD�6|C6D�D�:����8�?S̼�Q�?�,��+����?Q�y<�T]�~������D�6|C6D�D�:����8���n��M|?}�5?�<���=�q��U?~��=���D�+MC�e�D��0���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8������?Q���N�8�����>1�]�|b4��Z�	ݜ��yD�����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��N������&?�=����Q�z>1�]�|b4��Z�d���!Z�DW����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8����������������������������������������8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W���� 	 88�?x< >zMY    ���4�k�?�  >zMY�x< 4��ZC�c\B���    ���8��K�[�MGp?z��	�8�Q��>zMY�x< 4��Z������D2����8��a���c���Ԋ'>��=����h�>zMY�x< 4��Z@�@?����&����8�>��`�wq����B�a��c���Ԋ(>ʤ�>�c�h��Dl�,Cn�D�P����8�?iPB=�}�>����ʤȾ�x?h��=� ��}Sr����Dl�,Cn�D�P����8�<�������?~�?~NR=���7?��! ?}Sq=���De9C��@D�W����8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��K�[�MGo?z��	�8�Q��>zMY�x< 4��Z�OF��Q �C�_{���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8���������������������������������������� 	 88�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8��a��c���Ԋ(>��=����h�>zMY�x< 4��Z������D2����8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8�?�              ?�              ?�              ���8����������������������������������������8����������������������������������������8�����������������������������������������$DCSS_JPC 2������Q ( D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �$DCSS_JSC 2������Q ( @BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                              =���BS HALT                                               =���BS HALT                                               =���BS HALT                                 	              =����                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �                                                            �$DCSS_MODEL 2������Q x�                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �                           
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                              �$DCSS_PSTAT ������Q       (  (     ����                                                                                    ������������                  �������������$DCSS_SETUP 	������QB�                B�          �$DCSS_T1SC 2
������Q      Cz      Cz      Cz      Cz      Cz      Cz      Cz      Cz  �$DCSS_TCP R������Q � 
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                   
 D�                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �                                                                  �$DCSS_TCPMAP  ������Q @                            	   
                                                                      !   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @�$DCSS_TUIRO 2������Q �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �$DCSS_TUIZN 2������Q 	 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �$DCSS_UFRM R������Q � 	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                       	 8�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      