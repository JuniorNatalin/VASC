A��*SYSTEM*   V8.2306       4/24/2014 A 
  *SYSTEM* *SYSTEM*  
�WVAMP_T   $X1  $X2  $Y1   L�WVAMPFC_T   $AMP_ENB  $DT  �WV_RAMP_T   $ENABLED  $SCHD_NUM   ��WVCFG_T � $GROUP_NUM  $WV_ACCEL1  $WV_ACCEL2  $MAX_FREQ  $MAX_AMPL  $MAX_DWELL  $DEBUG  $MAXPREWS  $DOUT_NUM  $DOUT_PULSE  $DOUT_SHIFT  $DOUT_TYPE  $USE_AEFRAME  $GDO_NUM   $GDO_PULSE   $GDO_SHIFT   $GDO_TYPE   $WEAVE_TSK   $WV_TSK_GP   $SUPPORT_CF  $CNVT_DONE  $RAMP_ENB  $RAMP_GRP 2 $MAX_NUM_SCH  $ACCTIME1_GP   $ACCTIME2_GP   $EXTACC1_GP   $EXTACC2_GP   $MODE_SW  $COMP_SWITCH  �WVPHASE_T  4 $WVECT  $DWELL  $TERMTYPE  $DOUT  $PEAK  �WVPAT_T  \ $WVPAT_ID  $PAT_NAME $USE_START  $NUM_PHASE  $START_PHASE $WEAVE_CYCLE 2 
 ��WVSTATE_T   $CUR_REL_VEC    P�WVWPR_T  � 
$CENTER_RISE  $RADIUS  $WV_AXIS  $WV_FRAME  $AZIMUTH  $ELEVATION  $WV_BLEND  $CONTINUOUS  $DWELL_TYPE  $EXACT_SPEED  ��WVSCHD_T  H $FREQUENCY  $AMPLITUDE  $DWELL_RIGHT  $DWELL_LEFT  $L_ANGLE  �OTF_WV_T 	�  $OTF_ENABLE  $GET_AMP  $RAMP  $OTF_WVSCH $ORG_WVSCH $FBK_WVSCH $STEP_AMPL  $STEP_FREQ  $STEP_LDWL  $STEP_RDWL  $AMPL_H  $AMPL_L  $FREQ_H  $FREQ_L  $DWL_H  $DWL_L  $CHG_AMPL  $CHG_FREQ  $CHG_LDWL  $CHG_RDWL  $INC_AMPL  $INC_FREQ  $INC_LDWL  $INC_RDWL  $FBK_AMP  $CYC_ST_TK  $COM_ST_TK  $CYC_NUM  $DWL_SYM  $CHANGED  $UPDATE  $DEBUG  �$$CLASS  ������       �$WVAMP 2�������     ?   @�  ?      ���������   ���������   ���������   ���������   ���������   ���������   ����������$WVAMPTYP 2 �������  ?   @�  ?��u?   @�  @O�?   @�  ?   ?   @�  ?   ?   @�  ?   �$WVCFG �������      `   `   
   2  �           =���                                              =���=���=���=���=���=���=���=���                                                              ��������������������������������                                                                                                                 
    ,   }   }   }   `   `   `   `     �   }   }   }   `   `   `   `     `   `   `   `   `   `   `   `     `   `   `   `   `   `   `   `       �$WVPAT 2������� 
T   SINE                        ��                   
     ��  ?�    '                ?�  ��                    ?�  ?�    '                ��  ��                ������������������������������������������������������������������������������������������������������������������������������   FIGURE 8                                          
 ?   ��                      ��                          ?   ?�                      ?   ?�                      ��                          ?   ��                      ������������������������������������������������������������������������������������   CIRCLE              ?                            
     ?�                  �����                      ���    ��                  ���    ��                  ���?�                      ���    ?�                  ���������������������������������������������������������������������������������������   SIN 2                   ��        '             
     @         '              �         '          ������������������������������������������������������������������������������������������������������������������������������������������������������������������������   L                                                 
     �5)�5)  '                ?5)?5)                  ?5)�5)  '                �5)?5)              ������������������������������������������������������������������������������������������������������������������������������   Triangle                                          
     ��        '            ?�  ?�                      ��  ?�        '                ��                                                                                                                                                                                                 SINE                                              
     ��        '                ?�                          ?�        '                ��                                                                                                                                                                                                 SINE                                              
     ��        '                ?�                          ?�        '                ��                                                                                                                                                                                              ����              ��������������������������� 
 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������              ��������������������������� 
 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$WVSCHEXTENB         �   �$WVSTATE 2�������  �������������������������������������������������������������������������$WVWPR �������                                    �$WV_OTF 	�������            ?�  @�  =���=���    ?�  @�  =���=���    ?�  @�  =���=���    ?   ?   =���=���A�  =���A�  =���@�  <#�
                                                                �$WV_OTF_GP 2	�������  �            ?�  @�  =���=���    ?�  @�  =���=���    ?�  @�  =���=���    ?   ?   =���=���A�  =���A�  =���@�  <#�
                                                                