��   �*�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�NIO_AN_T�   L $�A* DR  �7SHIFT>V�ALID>I:I�E	IR�&CFG�.� �$V�ERSION �$COMME�NJ �USTOM� @ �2�DE_V_ENB> � �N�TMP�ST�ART_MODE~�NUM_LSJ��� �CHG_�DIG_PR�P�S_MAX���$� ;OP?] MKW>We�STr� ?I_OFS6O�] ��@q�����D<� KDV- KHO�L!�DH*ACT?_INDEX�c!�OPC�o!Kf*Kt)INIT�o �NNOT_NAM�� �$ORDE�= � �#HWl#�"R�EV�(SW1�*2r�*3#� SLO$�� VV3D 8IN��CP16XX_W&C51�D4��C53Y9PKX:PK~�SEARCH�� CHK�TP_�WA� c G�;M�AIN� Q>�2P�ARAM�7EXEyC6�R1SH2�S �HENABL�EpO^#SG_U}O�WD_TI� �;@ C� � P_DoEBUGPBSC,�?CS!DEFAUL�TPB�5�CAPD}U�PWRCLH<�1�KN_IO�A�K��!C�H�F�CFLA�G^#U!P�PWOFF_ALA� �BR� c"DBW@V��0�C.W�C�"2SY�;T[IO� �BOARD_S�!9B�T6�OP�YABD �XP�XMIS�U��W�ALM�Z�W��@`�U>A�Z� �YSM�VH�R� �XDc!iT�[�WmNOP fREAD�0�TS�T�D�fQ�1�j2�j3�UUP�DAT��0RC_�FIN@��aSI�Z�gJD�e>B�eDE��uPTH�fGR�OU��cOUJULONG�!Nt�!NtT1Nt4Kw5Kw6Kw�7Kw8KsBYTE �C�r�C�r1�tvq�t �q�t�q�t�q�t�q�tM9�w10��x1�x�1�x ��x1�x1��x1�x1�2����2. (d�f F)@�DI)0�ELTA#���	O�PT��W܆IOR_TRAN��ڄ�!RST�0��a��RESE�^PLI��1�S�"�INT#VL`L&X��O�!d�HO!$@ڀ�`@�ڀ�`@�U@RT�#���#��3�� vq���q���q���q�� �q���������(� ���@��ҙX���8p���FW_���1� 5 ��Wa�cN�CFIR�P@� ��&DB. �{ �
BASE�V) � UsI��� vs��vs�료s���s�/�뢈���Y�T��6��~�y�Pb{���o � �RE�@p��>A!5LAYw���bt��}ADD �@�W��W�t3W� �T�5\�6\�7\�8���IA� �� ���!$CNaT��uP�6��RI����PROC�`���` ���`�źB�D ����0�#�5Ϙ||�ǘ� A� �"X0���վ ��TYP������IP: < �����MAS�0��;pT�� ���QMSC�=�� �PrP>�Q�")�چ� O��"�D�!tF�UNK� �F��EXIl�C*`BUSY~���6*`�5��P� �槃@ B� U�Pr�F��FWV��SN��H���X1�`��� ��OCEX� A���� MAC��ML{FB��F_IP-����F_GW3�R3_1&U�U��SàCOU� �Ap�P1�� �� >AX3>A�>At3>Ay� >A��>A��>A��>A���� O�B��O���Z� ��e���p���{����s���s�USX3Oj� Pt3O��O��O��PO��O�� ��L��� � $PA�TH_XDЀA ����	c�� 	c� (u#���N��E�� ����$DOWN�LOA�9@�ARA�܀�#M�" ��L���l u����ً������S�NU�K_��&�K8! B�OPER@�8�A��CHE��J!��D$	bhS%�#	cB:�	2A'CPYA%��#LO� ^&�11A'�1�O(SE�R&��A'P ���'��B!��&�&t1�(��eB�K$�@0BUP� Y�5R e&.6�2�'�#7�!7 �"���)���)���)����#�a_BT'#�2DTV�5���3�d�5�6 B!���C�5�C�5�s�5 �s�"�8��D��D�� ,D��@�'�RvG5P���BADb@�WNGsGS�G$�TIN:`N�EAFE��@_��&��LD�9I�A=���P���P��SERVLI,�(�h!o���{���#CM:WSVFZLOIW	b��fW��NR���'IO5��V곐�в�pU�U��"�~dMOn�b$H!CM� �S��b�@t�NY�e a#c�tet�.f+�D&d�CLzf0�_+���ID _� [�lge�lg o�lg��lg��lg��ްYNC_�vc�e�c �bsf�e�k�c�e�c�e��c�e�cHp� L�1v��C!C! �s!�s!�s!�s! �s!�s!�Nr�Nr|Rw(�CLASS�`[����ve�������L� 	 � }ΪENABL����ES��+PENG�THJ>��_�UB09������DA7�S��]�ϠR�ERRDE�AC�I#�NDEX��3p���VPaQ�b�h��IM0x
�� $��H�"��L"��ET���V�񇠉Hٰ�bR5�0�B�F�"I#�����R_�N`P QIALB�$R7�0<Q1���$VMA��M.TSIMS��El���" ���AƠ � 
Ϊ9���>�㤽��PU%�摝��� ��]�_�4�������WRKxH 1v;v��	����`0�"�\�TP_DEBUG�"гO��_�PWO*0"�!W � �a�Ns��������ɥ�OM����U�BYT�����$S_�SYSY����U�g��yϋϝ��$�s  �����Y�a� N��#AN 2� ��N� M�� ������$��Խ�ǲ��ǲI�ǲ
-�ǲEςǲ]�ǲȰwϽ�$��ǲ��ǲ��ǲH���Ͻ���ǲߒǲ�ǲ 5�ǲ"$M�ǲ$e�ǲ&}�ǲI(��ǲ*��ǲ,��ǲ.��ǲ0�߂��"�CFG ���V820P02 131028�����O���P�־�	 ��� �~� �ś�@������X�� X��FANUC Ro�bot Cont�rollerC��A05B-260�0-J93 ��V�|�� � � !�Y� ��Y�dzm������� �����U��, ���e���f��mc:pniot?rc.txtX��ı��X�����{��2 "�L�B�&��N�C�y����װ����\) �b�젴� 2�� h�CP1604� DAP V2.�6i�L�!"�X�#$"�p�%"���'"���)5"��7"�)"� ��1m�L�� "�(M������0����16���+=Oaya����
�XX{i���/"/ �O/�/�/�/�/? %?7?I?[???�?�? �?�?������C��?O(O�?I���G ��!� .1�.��tM�1� �?�T۟TtO7O�ID���� �k�jltvl411�550r01rs--kux�O	__-_?_Q_���V_z_�_��_�_�_�__WS7-PC�_oo,o>o Poboe_�o�o�o�o�o��o�j!172.�26.29.20<hO�c255.&uB�bw�V"�=Z ~�c����� ���&��m6�Z�C� ~�m�����Ə���ُ8�V u�) ��!�Y�k�}���𡟳�ş�=L ���AMC:PC?ST_1.X� ���+�AUD1:�PN2610.FWL .3.9I�ql+�i����X�d d������� ����ʯܯ� ��jo 6�H�Z�l�~�����7��FR:S7PR�J�ֿ�9���\�fw_image.fwW�!�.�U��g�y��� ,X����h�|��@n[ ���H��@���C���� x��e�e�g����EEE������(��z (g��^!!����7�d��r	y���ST 2	d�J��D{?5�?����˓�p?����א������E���H�!�� K�5��Y��*�����AJ^����������!�"� �U����*���=�������<1������ ������� $6F�Hl~M� ������2 DV%z�[�� ���
//�@/R/ d/3/�/�/i/�/�/�/ �/??*?�/N?`?r? A?�?�?�?�?�?�?�? O&O8OO\OnO�OOO �O�O�O�O�O�O�O_ 4_F__j_|_�_]_�_ �_�_�_�_oo�_Bo To#oxo�o�oko�o�o �o�o,�oPb 1t��y��� ��(�:�	�^�p��� Q�������܏� �Ϗ $�6�H��l�~���_� ��Ɵ��؟���ݟ2� D�V�%�z�����m�¯ ԯ毵�
���@�R� d�3�������{�п� ��ÿ�*���<�`�r� AϖϨϺω������ ��&�8�J��n߀�O� �߶��ߗ�������� 4�F�X�'�|��]�� �����������B� T�f�5�������}��� ����,��Pb tC������ �(:	^p� Q����� // �6/H//l/~/�/_/ �/�/�/�/�/? ?�/ D?V?%?h?�?�?m?�? �?�?�?
OO.O�?RO dOvOEO�O�O{O�O�O �O�O_*_<__`_r_ �_S_�_�_�_�_�_o �_&o8oJoono�o�o ao�o�o�o�o�o�o 4FX'|��o �������0� T�f�5�������}�ҏ ���ŏ�,�>��b� t�C������������ �ӟ(�:�L��p��� Q�����ʯ��� �� �6�H�Z�)�~����� q�ƿؿ����� �� D�V�h�7όϞϰ�� ���ϵ����.���R� d�v�Eߚ߬߾ߍ��� �����*�<��`�r� ��S��������� ���8�J��\����� a�����������" ��FXj9��o ����0� TfxG��}� ���/,/>//b/ t/�/U/�/�/�/�/�/ ?�/(?:?L??p?�? �?c?�?�?�?�? OO �?$OHOZO)O~O�O�O qO�O�O�O�O_ _2_ _V_h_7_�_�_�__ �_�_�_�_o.o@oo dovoEo�o�o�o�o�o �o�o*<Nr ��e����� ��8�J�\�+����� ��s�ȏڏ����"� �F�X�j�9������� ��֟���ɟ�0��� T�f�x�G��������� ����ׯ,�>��P� t���U�����ο��� ���:�L�^�-ς� ��cϸ����ϫ� �� $���H�Z�l�;ߐߢ� qߴ����߹�� �2� �V�h�z�I����� ���������.�@�� d�v���W��������� ����<Nr ��e���� &�J\+�� �s����/"/ 4//X/j/9/|/�/�/ �/�/�/�/�/?0?B? ?f?x?�?Y?�?�?�? �?�?O�?,O>OPOO tO�O�OgO�O�O�O�O __�O:_L_^_-_�_ �_�_u_�_�_�_�_o $o�_HoZolo;o�o�o �o�o�o�o�o�o 2 DhzI��� ���
��.�@�R� !�v���W�����Џ�� ����<�N�`�/� ����e���̟ޟ��� �&���J�\�n�=��� ������گ쯻��"� 4��X�j�|�K����� Ŀ�����ɿ�0�B� �f�xϊ�YϮ����� ��������>�P�� t߆ߘ�g߼����߯� ��(���L�^�-�p� ���u��������� $�6��Z�l�~�M��� ������������ 2 Dhz�[�� ���
�.@R�!v��e�$P�NIO_IM0 �
�����N�k�� V�A05B-260�0-J930e�F1732681 ��k���LST 2	�DXn;*�?�e�F'P_$g|/K#�i$�Z/(l/�/"H� �$� !�/�/�/�"�!�/?�=J�(*?<?N??��y4ʞ/|?�?L"�`�8�#�?OC*�$p�1)?OO �.H m?KO�O�O]�O�O�O �O_0_B__f_x_�_ Y_�_�_�_�_�_o�_ ,o>oPooto�o�ogo �o�o�o�o�o( L^-���u� ����$�6��Z� l�;���������؏� ��ˏ �2�D��h�z� I����������
� ٟ.�@�R�!�v����� i���Я������� <�N�`�/�������w� ̿޿����&���J� \�n�=ϒϤ϶υ��� ������"�4��X�j� |�Kߠ߲��ߓ����� ���0�B��T�x�� Y����������� ��>�P�b�1�����g� ��������(�� L^p?��u� ���$6Z l~M����� �� /2/D//h/z/ �/[/�/�/�/�/�/
? �/?@?R?!?v?�?�? i?�?�?�?�?OO*O �?NO`O/O�O�O�OwO �O�O�O�O_&_8__ \_n_=_�_�_�_�_�_ �_�_�_"o4oFoojo |o�o]o�o�o�o�o�o �o0BT#x� �k������ �>�P�b�1������� y�Ώ������(��� L�^�p�?��������� ܟ� �ϟ$�6��H� l�~�M�����Ư��� ���ݯ2�D�V�%�z� ��[���¿Կ����
� ��@�R�d�3ψϚ� iϬ����ϱ���*� ��N�`�r�Aߖߨߺ� �����߿��&�8�� \�n��O������ �������4�F��j� |���]����������� ��BT#x� �k���� ,�Pb1t�� y����/(/:/ 	/^/p/�/Q/�/�/�/ �/�/ ?�/$?6?H?? l?~?�?_?�?�?�?�? �?O�?2ODOVO%OzO �O�OmO�O�O�O�O
_ _�O@_R_d_3_�_�_ �_{_�_�_�_�_o*o �_<o`oroAo�o�o�o �o�o�o�o&8J n�O���� ����4�F�X�'� |���]���ď֏���� ���B�T�f�5��� ����}�ҟ䟳��� ,���P�b�t�C����� ���������(�:� 	�^�p���Q�����ʿ ��� ���6�H�� l�~ϐ�_ϴ����ϧ� ��� ���D�V�%�h� �ߞ�m������ߵ�
� �.���R�d�v�E�� ��{����������*� <��`�r���S����� ��������&8J n��a��� ���4FX' |��o���� //�0/T/f/5/�/ �/�/}/�/�/�/�/? ,?>??b?t?C?�?�? �?�?�?�?O�?(O:O LOOpO�OQO�O�O�O �O�O __�O6_H_Z_ )_~_�_�_q_�_�_�_ �_o o�_DoVoho7o �o�o�oo�o�o�o�o .�oRdvE� �������*� <��`�r���S����� ̏�������8�J� �\�����a���ȟڟ �����"��F�X�j� 9�����o�į֯请� ��0���T�f�x�G� ����}������ſ� ,�>��b�tφ�UϪ� ���ϝ������(�:� L��p߂ߔ�c߸��� �߫� ����$�H�Z� )�~���q������� ��� �2��V�h�7� ��������������� .@dvE� ������* <Nr��e� ���//�8/J/ \/+/�/�/�/s/�/�/ �/�/?"?�/F?X?j? 9?�?�?�?�?�?�?�? �?O0O�?TOfOxOGO �O�O�O�O�O�O_�O ,_>__P_t_�_U_�_��_�_�_�_oo�R��$PNIO_MO�D 2����;aN� � @DAP OV2.6o�Phd�j`ka�_SAF�E 8 BYTE�zohchd{oS32�o�Vhd7hc$�fka �o~hdUa �d�b�as^p�_ �������� $�6�	�Z�l�?����� ����؏ꏽ�� �2� �V�h�;�z������� ԟ���˟�.��R��d�v�+gSTM  =;eNja+q ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x����O_WRK �;i ���_j|�bC���X�� �