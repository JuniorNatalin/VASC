��   &�A��*SYST�EM*��V8.2�306 4/2�
 014 A �	  ���C�ELLSET_T�   w$�GI_STYSEL_P 7_T  7ISAO:iRibDi�TRA�R��I_INI; ���t�bU9ARTaRSRPNS1Q�2345*678Q
�TROBQACKSNO��) �7�E�S�a@�o�z2 U3 4 5 6 �7 8awn&GINm'D�&��)%� �)4%��)P%��)l%3SN�{(OU��!|7� OPTNA�73�73.:B<;}a6�.:C<;CK;CaI?_DECSNA�38R�3�TRY1���4��4�PTHC�N�8D�D�INCYC@HG�KD�?TASKOK�{D �{D�7:�E�U:�C h6�E�J�6�C�6U�J��6O�;0U��:IAT�L0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T��T�@REQ�d��drG�:Mf�GJO_HFAUL�Xd�dvgALE� �g�c�g�cvgE� �H�dvg�NDBR�H�dgR�GAB�Xtb ��CLMLIy@�   $�TYPESIND�EXS�$$CL�ASS  ����lq������$'61ION  �����q}t+ UP0 lu�q�Style�-Auswahl�	  ��r�t A�nf./Echo��s�zck����ystarten���t"�1�C�XR�d�  
����U���������q�������q�r�s�Option B�it A �ʎB�܏҆C���tcod�e�w�tTryou?tmodus�w��Bahnseg. weiter��In ZyklI���Aufg OK��Manuel� Ѐ.�qA����B4����Cܜ. �t�q��yRoboh�ve�rria�� � i�n Isolat�e��{���\�ment�w�t\��pd��>@�-StatI���	MH Faul�t:����Aler|ϯ��#  ����	�}p@r 1�z �.��:�L�
�; L�E_COMNT �?�y�    ��Ɔ������ʿܿ�  ��$�6�I�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ�@����������r�U}������   r�E�NAB  �� ��W�i�{�����r�MENU �yt�NAME ?%��(%$*���&��p �M�8�q�\�x����� ����������7" 4FXj|��� ����WB {f������ �//A/,/H/P/b/ t/�/�/�/�/�/?�/ ??(?:?L?�?p?�? �?�?�?�?�=