��   ɋ�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�CSS_CPC_�T   � �$COMMENT� $ENA�BLE  $�MODJGRP_�NUMKL\ � $UFRM�\] _VTX �M �   $Y��Z1K $Z2��STOP_TY}PKDSBIO��IDXKENBL?_CALMD�&}S. � 8�J\TC�u
SPD_LI_����COL�&Y0 � � !CHG�_SIZ$A�P7ECDIS � � �7�C�����Jp 	�J �� ��"��$�'"_SEs�xSTAT/� D $FP_�BASE �$LINK`$!��j&_Vs.Hs# � �&J- ���ZAXS\UPR:LW�'CU��  �$� | 
�/�/�/4�??j&ELE�M/ T $1Uc c1j"NO�7�0�a3UTOOi�2H�A�4�� $DA{TA"  x&e0   @P:�0� 2 
&PNP% ��P!U*.n   oFSyCjHrB� zB(�F�D(�1�R5C�DROBOT��H�CQBo�E�F$CUR_"�B<4�SETU�	 l|� �P_MGN�INP_ASS�  @�� �3�8"7GP� U�>VhSP!��4T1�
@B\8�8�T= �0 P�+ Kec1V�RFY�8�T$5&1ȕ ��W��1$�R�UPH/ ([ �#A�#A�#A�3tBOX/ 8�0�����`bto%cԅTUIR�0  ,[ �62`�ERa02 $�k` �a_S��b��fZN/� 0 [9&0� LarZ_� �_� 8tu0  @�A�Y�v	�on�$$�CL,P  �����q��Q��Q��$' 2 �u�Q   �(�q���b0�p�}�p��~�4�F� ��m������Ǐ ُL�������E��� i�{���$�6�� Z�����A���Ɵ؟ ��������2��V�h� z�+���O�a�ԯ���� 
�@�Ϳ����v�'� �����п^ϓϥ�� ��<�N���r��5�G� ��k����ϡ������ ��\��ߒ�C��g� y��ߊ��"�4���X� 	����?�������� �����0���T�f�x� )��M_����� �>�t%� ��m\��� :L�p�3/E/� i/��q//�/�/�/ Z/?~/�/A?�/e?w? �?�/�? ?2?�?V?O O�?*OOO�?�?�O�? �O�O.O�OROdOvO'_ �OK_]_�O�_�O__ �_<_�_�_r_#o�_�_ �_ko�_�o�oo�o8o Jo�o�o1C�og �o�o"���X 	�|���O�u��� ����0��T��� )���M���ҏ������ ��,�ʟ�b�t�%��� I�[�Ο����ǯ :����p�!��������i�ܯ������$D�CSS_CSC �2I�ɱ?Q  D��� @���&���J�\�n� =ϒϤ϶υ������� ��"�4��X�j�|�K� �߲��ߓ�������� 0�B��f�x��Y�� �����������>� P�b�1�����g������������GRP ;2ɻ ��	��cN�r�� ����;& Kq\����� �/�%//I/4/m/ X/j/�/�/�/�/�/�/ ?�/3??W?B?{?f? �?�?�?�?�?�?�?O OAO,OeOPO�O�O�O |O�O�O�O�O___ O_:_s_�_T_f_�_�_ �_�_o�_'oo7o]o oo>o�o~o�o�o�o�o��o�o5
ST�AT 2ɹY��,8�?z��ͽ�g~�=J�-��f�xP��>w��Jz���liֿs����9�-�N���D�K�ɱ,p8~xq��wz����4��Z��T��?�p�q6�p�q����Ü�ɱxq6�&r�>�\�?b	M6�J�q���p�y:���C@�
DmKD�v�8��?��?�Y��q������ �6j���0��-�:���C��]D���u�>T�}?� �?T\^6v�0��H��zg��=�[>4�1��.10�Ahf�D�H�u������w{^>}��$?zg���Q�4�>Jz��>li�?s�؄�z��́ɵ� �ɵ�J�\�:����� �y�q����Ȇş� ٟ�%��!�3�E�W� y�{�����ٯ�v��� d��H�Z�8�~����� 䯺���ƿ�ڿ��&� �2�\�F�hϒ�|ώ� �ϲ�p�
����@�R��0�v߈�f�Ѐɽ��fY؀���lG��xQ0>wl�耧�lb��s��E�9��N��o�p&�z��{��&�i�v���q��t��~�JS>��[��p�6���$�!���:�΀�C@�����v��<�?�g?Y��4�􈜵 ��6��z\��Y�;1�fC���wT��X��?��?T]H6�&�\��t�hx��=��U���������Aj�D�G�Z���*���>}������K���尀�>lb�?s�D��߸��� l�>�P�.�t���d��� ������������ (R<N�r�� �����6H�� l~\����� �/�/2/4/F/ h/�/|/�/�/�/�/�/ $.?@?�d?v?T?�? �?�?���������� �&�8�J�\�n��� ����������?�?"� �?n_�?^_�_�_�_�_ �_�?o�/"oLo6o Xo�olo�o�o�o�o�o �o�o$�_fxV ������_8� �D�.�P�z�d�v� ������ΏЏ��.� �^�p��������ʟ ܟ�?,_>_�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__��R_ ��������Կ���
� ��<�F��R�|�f� �ϲϜϾ�������� �*�T�>�ϖ�迆� ���߼���.�h�>� D�J�t�^����� ������� ��L�6� �ߎ���~��������� ��\�n�,�>�P�b� t���������ί�� ��(�:�$6H�� �����/�(/:/  �J�d/n�`/�/�/�/ �/�/�/�/??$?N? 8?Z?�?v��?�?/�? �?�?O2OL/^/�?nO t?zO�O�O�O�O�O�O _�O_F_0_R_|_f_ DO�_O�_�_o�_*o <oz��\n�� ������" lFXjTofoxoo ���"�4��X�j� PO�_���_��ʏ��Ə  ����� �2�T�~� h������_���H�� ,�
�P�b�|�����ʟ ���������
���� @�*�L�v�`�����ҟ ܿ�@���$��4�Z� 8Ϫ���o�o�o�o �o�o�o
.@R dv��߄ϖ��J� �.��R�d�B��� ������������ 0��<�f�P�b����� ������z�&J \:��������� ����($F HZ|���� //pB/T/2/x/�/ t����ߪϼ������� ��(�:�L�^�p߂� �ߦ߸��ߴ/�/ �/ LO�/\O�O`OrO�O�O ���O� _*__6_ `_J_l_�_�_�_�_�_ �_o�_�ODoVo4ozo �ojo�o�o�Oo�o�_ �o".XBd� x�������o <�N�,�r���b�������e�$DCSS_�JPC 2�e�Q ( D��%��$�6�H� �l�~���_���Ɵ�� �����ݟ2�D�V�%� z�����m�¯ԯ毵� 
�����R�d�3��� ����{�п���ÿ� *����`�r�AϖϨ� �ω��������&�8� J��n߀�O�a߶��� ���������4�F�X� '�|��]�o������ ������B�T�f�5� ������}��������� ,��PbtC� �������( :	^p�Q�� ��� //�6/H/ /)/~/�/_/�/�/�/ �/�/? ?�/D?V?%?�7?#�؅S��@�BS HALqT�?u5u?  )�=��ʹ?�?�4!�?�?O�6 O2ODO�6`OrO�O�6�A�O�O�O�3�O�OC_B�6 _2_�_�6`_Hr_�_�6	�_�P��_ ox?$��_Eoo*o{o No�oro�o�o�o�o�o �o�oA&wJ\ n������� =��a�4���X�j��� ��ɏ���֏�9�� �0���T�f������� ����ҟ�"�G��,� }�P���t�ů������ ί	��C��(�y�L� ^�p���������ʿܿ �?��$�bχ�Z�l� �ϐ��ϴ������;���I�2߃�Vߊ?_MODEL 2�;�xt�i�
 <*m�c�:�H�J"� ���X�/�A�S�e�w� ������������ �+�=���a�s����� ����������g�P�� +�o���� ����L#5� Yk}��� /� �6///1/C/U/g/ =�/a�/�/?�/�/ D??-???�?c?u?�? �?�?�?�?�?�?@OO )OvOMO_O�O�O�O�O �O�O�O�/�/�/__ �_�Om__�_�_�_o �_�_8oo!o3oEoWo io�o�o�o�o�o�o�o �ojAS�;_ M_{��u��� �+�x�O�a������� ����͏ߏ,���b� 9�K�]�o��������� ɟ�����p�� Y�k��������ůׯ $�����l�C�U��� y���ؿ����ӿ ��� 	�V�-�?ό�'�9�K� yϋ�a�����.��� d�;�M�_�q߃ߕ��� ���������%�7� I��m�������� ��&��������E�W� ��{������������� ��X/A�ew ������B +=��7�ew ���/�/P/'/ 9/K/�/o/�/�/�/�/ ?�/�/�/L?#?5?�? Y?k?�?�?�?�?�O ��?�?ZO1OCO�OgO yO�O�O�O�O_�O�O D__-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o�?�o#OQoco�o�o �o�o�o%7 �[m����� ��8��!�n�E�W� i�{�����uo���oǏ ُF��/�|�S�e�w� ğ������џ�0�� �+�x�O�a������� 䯻�ͯ߯,���� ���=�O���7����� ɿۿ�:��#�p�G� Y�k�}Ϗϡ������� $�����1�C�Uߢ� yߋ���s�������2� ���-�?�Q�c��� ������������� d�;�M���q������� ������N���� );�#���� �&�\3EW �{����/� �/X///A/�/e/w/ �/_q��/�/�/? ?f?=?O?�?s?�?�? �?�?�?O�?OPO'O 9OKO]OoO�O�O�O�O�_�O�O�O�$�$D�CSS_PSTA�T ����cQQ   g t_�Z r_ (�_�_�WkPkP�_n�_ l c�dP��P;_4oFo�)�"ocUcUdovoTTSE�TUP 	cYB�&T�#�!�dOYT1SC 2
�j`�!Cz�#|/}�eCP R�l�� DSoz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ��.h%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛ�� ���������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�����}� �������������� 1CUgy�� �����	- ?Qcu�������Z�D�/*/</ �/`/r/�/S/�/�/�/ �/�/??�/8?J?? [?�?�?a?�?�?�?�? �?O"O�?FOXOjO9O �O�O/}O�O�OoO_ _0_�OT_f_x_G_�_ �_�_�_�_�_�_o,o >ooboto�oUo�o�o �o�o�o�o:L �O)����� � ��$��H�Z�l� ;�����q���؏ꏹ� � �2��V�h�z�I� ���������_՟ .�@�ǟd�v���W��� ��Я�������<� N��_�����e���̿ ޿����&���J�\��n�=ϒϤ�s��$D�CSS_TCPM�AP  ������Q W@ ~�~�~��~���~�~��~�~�	g�  �~�~�~�~��~�~�~�~��~�~�~�~�R~�~�~�~�~�U~�~�~�~�U ~�!~�"~�#~�U$~�%~�&~�'~�U(~�)~�*~�+~�U,~�-~�.~�/~�U0~�1~�2~�3~�U4~�5~�6~�7~�U8~�9~�:~�;~�U<~�=~�>~�?~��@��UIRO 2]�����$� �"�4�F�X�j�|�� �������������0�B�T�}��}�� ������������ 1CUgy��� ��^�����-? Qcu����� ��//)/;/M/_/ ��/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?�?�?�?v/O���UIZN 2.��	 �����PO bOtOy�KO�O�O�O�O �O�O_�O0_B_T__ x_�_�_k_�_�_�_�_ �_o,o�_Poboto�o Io�o�o�o�o�o �o:L^-��� i�����$�6� �Z�l�~�M�����Ə ؏�����ݏ2�D�V��O��UFRM R�����џ��� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߒ��� ������������/� A�S�e�w����� ��������+�=�O� a�s��ߗ��������� ��'9K]o ���������#5GYk���x������ //�B/T///x/�/ e/�/�/�/�/�/�/? ,??P?b?y��?�? I?�?�?�?OO�?:O LO'OpO�O]O�O�O�O �O�O�O�O$_6__Z_ l_�?�_�_A_�_�_�_ �_o�_2oDoohozo Uo�o�o�o�o�o�o�o .	Rd{_�� 9������� <�N�)�r���_����� ��ޏ��ˏ�&��J� \�sw