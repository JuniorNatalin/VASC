��   ��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�MC_CFG_T�   � $�'NUM_MSK�  $EXE�_TYPECME�M_OPTPN_�CNFCIF_C�Y:gSCN_T�IME E RESET_P�Do �LJ �HECK_�DSBLC $D�RA> ARGIN�CSTORJ  ݼ&DEV. �d 	7OC'H�AR�ADD�S�IZORACBS�LO[ODKIO>KOCCPYC&|l /  L ���h99IDX�C��&L. 7� 
�EQPLnHRAT�TRK�BUF| ��U�N_STATUS�CU��MAX�(I�-<�S�NP_PA�  �� � AN�NE�� OW CToION_�PU��   $B�AUD�NOIS�YmN�T1�#2��#3�$_PR�Ty4P' DATA��CQUEUE� P;TH[$MM_��%�&!RETRIES^CAUTO!R[���BG � �I?SP_INFd�<' CLIMI� B5AD_H C3H��# d6�#d6�#d6�#W1� ��#�4�#�4�#�4�" �`�$$CLA�SS  ��i��1�����i�FG0 �5���C�2��� B�d��C�3�  2:�7	@d $DZO ��WO�O{O�O�O�O�O �O�O__@_/_d_S_ �_w_�_�_�_�_�_�_ oo<o+o`oOo�oso �o�o�o�o�o�o 8'\K�o�� ������4�#� X�G�|�k�����ď�� �׏���0��T�C� x�g����������ӟ ���,��P�?�t�c� ���������ϯ�� (��L�;�p�_����� ����ܿ˿ ��$�� H�7�l�[ϐ�ϴϣ� �������� ��D�3� h�Wߌ�{߰ߟ����� ������@�/�d�S� ��w���������� ��<�+�`�O���s� ������������ 8'\K�o�� �����4# XG|k���� ��/�0//4,�3�IF 2CKP �DXD�G�%U�@@!�,�$T"A�)�$�,��$U�+A@<(*�!�()DY�(1H�%/0�&"<<�%<<�%<<�%	<;6EP�55S1'5F�(�(��1�!�!�;�"�!��<�� H@��8G��(,L�5,K
F\L#E��8K�4k10�'k5�@��4�A�ڜ4R�3�3*��4D�3�@C�F7@
C"H@DA�7�F�1U &_!_3_E_n_i_{_�_ �_�_�_�_�_�_oo FoAoSoeo�o�o�o�o �o�o�o�o+= fas����� ����>�9�K�]� ��������Ώɏۏ� ��#�5�^�Y�k�}��������şS/e"TY�PE 2o+ �(�3�!d�6�|蟮1�ڞ�0 L���ZAt����!��կ����b!SNP_PARAM o+"ΥϯƧ�A'� S� ̦�0[A�"�1l��1�!U&��)4�