��  IL�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���S�BR_T   �| 	$SVMT�R_ID $R�OBOT9$GRP_NUM<AXISQ6K 6�NFF3 _PA�RAMF	$�  ,$MD �SPD_LIT U�&2*� �� �s@p�$$�CLASS  ������ � ��$'  1 ���  T����R-2000i�B/210F���ACaiS�R30/3	 8�0A��
H1 DSP1-S1���	P01.05�,  	��  ��Pa�R���b��w���������
=�#�,r�9  ~���%����8� l� � ����?� %����(�� �����l��k��/  �3!���=������=���vG�����&��S � ���� �m��������ǣ�Z �I���yH!��j�����c9	`�B 0 ���� �� :?p��@  'bx�'/�/�/�/�/��3�/�/3 ?%?�7?��Z��3�!�������e���3@������� 
�'�#!>?�?�, )$62@2HZrl�� �8�D�֞��h�� ���  ������ 3��f��<�����wDӿ�7�D *#�  ����� O$� �O�������>'��2^ Q
��(T(�`/ r/�!@�/T_f_x_�_��/�_	?�_�_??Q? �3E�������N	5��5k
}���;w�/��
�?
k'�:�_Uo&���?�?6�3@�ROK��q��\�3�cDO���phOz@y�/ǫ/����D^4��դ@����Fw�4t0���K����@��� 6R$v\o����@K>(���	��9��ST(�_*_<_ ��)�;��__��_p� ����oˏݏ���s�po�`�12/41�S 4�5;4@4�o�m�z�e�q��f��2�"<C�p�d?�k0������ (H������ܕ@�� ��@�7A$A@������@��� ;$��'��D��0>!�]����VP���@�����  ��������s~"��y ���ɯۯ���Z�#��f(�M�_�q����������˿�b,�L�^�5@{�t�������8G�ݴ�Ɵؕ�
���!!�>��>�������5���>�Cd����������f�N�>x����`�������u߇ߙ߫� ���*�����)�;�0M�_�q����	�^�6@�r,�>��P� `�$l�~����ܑ�� =��LL��}�����* ��SD ���E�f����<��
�o�U�~�.@� R�d�-?Qc�߇ �ߘ�����);M�����<TqPPgu	u��o�� ���//,/>/P/ b/t/�/�/�/�/�/�/�/?<�?8?J?\? n?�?�?�?�?�?�?�? �3n`
O���pO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_"?�_�_o o 2oDoVohozo�o�o�;�  =�EX�TENDED A�XIS���q?aiS4/5����nAAH h� -ND���0.3����  �P���r  H��X�o������  {�'�9�~�5
�� ��� ��l� �ܑt�Ƃ������� ���c	`� 7 (���t Z�	�!�_�q�����������ӏ叀��	��-�?�Q�c��(OO|�>OPObO� ����*�<�N�`�r� ��������̯ޯ�� �&�8��_\�n����� ����ȿڿ�����? ����Yϴ�Ɵ�Ϡϲ� ����������0�B� T�f�xߊߜ߮����� ��@���,�>�P�b� t�������*�<� ��`�rτ�L�^�p��� ������������  $6HZl~�� ������ 2 DVhz����� �0�B�
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?� �?�?�?�?�?�?�?O O&O8O����O� ��O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oh?0oBo Tofoxo�o�o�o�o�o �o�oROdO�O�O�O t������� ��(�:�L�^�p��� ������ʏ&o� �� $�6�H�Z�l�~����� �o0"̟FXj2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���䏬���п� ����*�<�N�`ϼ� ������������ �&�8�J�\�n߀ߒ� �߶����������"� 4X�j�|���� ����������zό� 6������Ϝ������� ����,>Pb t������� N�(:L^p������&�  =��EXTEN�DED AXIS�h���aiS�4/5000 4�0Ak�H  D�SP -~�P0�0.39�� 	o�  o�Pm�} H�X�q������  �{n�C 9~��5
�� �p� �l�� l���tn�b��/�/�/��/
??.?e�c�	`� 7 �(�"t Z� �:?=�j��!>?�?0�?�?�?n��?�? OO'O9OKO]OoO�O�O�X�J��On��� ��_$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVoho�o�o �o�o�o�o�o
. @,��O�O��O�O� �����*�<�N� `�r���������̏ޏ ����po8�J�\�n� ��������ȟڟ��� Zl����|��� ����į֯����� 0�B�T�f�x������� ��ҿ.�����,�>� P�b�tφϘϪ��� *i!/%/7/I/[/m/ /�/�/�ߦ߸����� �� ��E?W?i?{?l� ~����?�������� � �2�D�V�h��O=� /���S�e�����	 -?Qcu��� ����); ߿Mq����� ��//%/���=/ �������/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?U O/OAOSOeOwO�O�O �O�O�O-/_/Q/�Ou/ �/�/a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�oO�o �o�o#5GYk }��O__�3_E_ ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c��ou����� ��ϟ����)�;� M���e����˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�}�E�W�i�{� �ϟϱ���������U� ��y�#ߝ������ߛ� �߿���������+� =�O�a�s����� ����;���'�9�K� ]�o����������E� 7� [�m�5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�����/ +�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO� mOO�O�O�O�O�O�O �O_!_}/�/�/K_�/ �/�/�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�ocO+ =Oas���� ��;_m___(��_�_ ]�o���������ɏۏ ����#�5�G�Y�k� }�������ş��� ��1�C�U�g�y��� ������/�A�S�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�q�͟�ϧϹ��� ������%�7�Iߥ� ׯɯs��������� ���!�3�E�W�i�{� ������������� �/���S�e�w����� ����������cߕ� ��P�߽߅��� ���'9K ]o������ 7��/#/5/G/Y/k/ }/�/�/�/�/!3�/ Wi{C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O� �O�O�O�O__)_;_ M___q_�/�/�/�_? '?9?oo%o7oIo[o moo�o�o�o�o�o�o �o!3EW�O{ �������� �/��_�_�_x��_�_ ����я�����+� =�O�a�s��������� ͟ߟ��_�9�K� ]�o���������ɯۯ �I�[�������k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ��������	�� -�?�Q�c�u߇ߙ��� '����=�O�a�)�;� M�_�q������� ������%�7�I�[� m���ϣ��������� ��!3EW���� �ߠ������ /ASew�� �����//+/ ��=/a/s/�/�/�/�/ �/�/�/??q�-? ����?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�OE/ __1_C_U_g_y_�_ �_�_�_?O?A?�_e? w?�?Qocouo�o�o�o �o�o�o�o); M_q���_� ����%�7�I�[� m���_o�_ȏ#o5o ���!�3�E�W�i�{� ������ß՟���� �/�A�S��e����� ����ѯ�����+� =�����U�Ϗ�󏻿 Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����m�5�G�Y�k� }ߏߡ߳�������E� w�i�����y�� �����������	�� -�?�Q�c�u������� ����+���); M_q����5� '��K�]�%7I[ m������ �/!/3/E/W/i/{/ ���/�/�/�/�/�/? ?/?A?S?e?��}? �	�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_�/ ]_o_�_�_�_�_�_�_ �_�_om?�?�?;o�? �?�?�o�o�o�o�o�o 1CUgy� ������S_� -�?�Q�c�u������� ��Ϗ+o]oOo�so�o M�_�q���������˟ ݟ���%�7�I�[� m���������ٯ� ���!�3�E�W�i�{� ��������1�C�� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a߽��ߗߩ߻� ��������'�9 ǿ��c�ݿ������ �����#�5�G�Y�k� }��������������� {�CUgy� ������S�� w�@���u��� ����//)/;/ M/_/q/�/�/�/�/�/ '�/??%?7?I?[? m??�?�?�?#�? GYk3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�/ �_�_�_�_�_oo+o =oOoao�?�?�?�oO O)O�o'9K ]o������ ���#�5�G��_k� }�������ŏ׏��� ��{o�o�oh��o�o ������ӟ���	�� -�?�Q�c�u������� ��ϯ��O��)�;� M�_�q���������˿ ݿ9�K���o�����[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱��������� �/�A�S�e�w��� �	ϳ�-�?�Q��+� =�O�a�s��������� ������'9K ]o�ߓ���� ��#5G���� ���������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? w-?Q?c?u?�?�?�? �?�?�?�?OasO ����O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_5? �_o!o3oEoWoio{o �o�o�oO?O1O�oUO gOyOASew�� �������+� =�O�a�s������_�� ͏ߏ���'�9�K� ]�o��o�o�o��% ����#�5�G�Y�k� }�������ůׯ��� ��1�C���U�y��� ������ӿ���	�� -ω���EϿ�џ㟫� ����������)�;� M�_�q߃ߕߧ߹��� �����]�%�7�I�[� m���������5� g�Y��}Ϗϡ�i�{� �������������� /ASew�� �����+ =Oas����%� ��;�M�/'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? �}?�?�?�?�?�?�? OO1OCOUO��mO ��/�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o�? Mo_oqo�o�o�o�o�o �o�o]O�O�O+�O �O�O������ ��!�3�E�W�i�{� ������ÏՏ�Co� �/�A�S�e�w����� ����M?�cu =�O�a�s��������� ͯ߯���'�9�K� ]�o������ɿۿ ����#�5�G�Y�k� }�ٟ럕��!�3��� ��1�C�U�g�yߋ� �߯���������	�� -�?�Qﭿu���� ����������)��� �ϩ�S������Ϲ��� ����%7I[ m������ �k�3EWi{ ������C�u� g�0/����e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?OO'O9OKO ]OoO�O�O�O//�O 7/I/[/#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�? �o�o�o�o�o�o	 -?Q�O�O�O{�O __����)�;� M�_�q���������ˏ ݏ���%�7��o[� m��������ǟٟ� ���k��X��� ������ïկ���� �/�A�S�e�w����� ����ѿ�?����+� =�O�a�sυϗϩϻ� ��)�;���_�q���K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }������������� ��1�C�U�g�y��� ��ϣ��/�A�	 -?Qcu��� ����); M_������ ��//%/7/���� ���/�����/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O gOAOSOeOwO�O�O �O�O�O�O�OQ/c/_ �/�/�/s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o%O �o�o#5GYk }���O/_!_�E_ W_i_1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u����o�� ��ϟ����)�;� M�_�������� ݯ���%�7�I�[� m��������ǿٿ� ���!�3Ϗ�E�i�{� �ϟϱ���������� �y���5߯���ӯ�� �߿���������+� =�O�a�s����� ������M��'�9�K� ]�o�����������%� W�I���m�ߑ�Yk }������� 1CUgy� ������	// -/?/Q/c/u/�/�� �/+=??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O �mO�O�O�O�O�O�O��O_!_3_E_�$�$SBR2 1�%�qP T0 '� �/�) �_�_ �_�_�_�_oo,o>o Poboto�o�o{_�_�o �o�o(:L^ p�����o�o�o  ��$�6�H�Z�l�~� ������Ə؏��� �2�D�V�h�z����� ��ԟ���
���� @�#�d�v��������� Я�����*�<�N� 1�r�U�������̿޿ ���&�8�J�\�n� ��c�L_���������� ��,�>�P�b�t߆� �ߪ߸ٚ�������� "�4�F�X�j�|���������� � ���#�5�G�Y�k�}� �������������� ��0BTfx�� �����, >��bt���� ���//(/:/L/ ^/p/T�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�/�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�?�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_o�O*o<o No`oro�o�o�o�o�o �o�o&
oo\ n������� ��"�4�F�X�<h� ������ď֏���� �0�B�T�f�x���n� ����ҟ�����,� >�P�b�t��������� ������)�;�M� _�q���������˿ݿ �"�$�6�H�Z�l� ~ϐϢϴ��������� � ߤ�D�V�h�zߌ� �߰���������
�� .�@�R�6�v���� ����������*�<� N�`�r���د������ ����'9K] o����j��� �"4FXj| ��������/ /0/B/T/f/x/�/�/ �/�/�/�/�/?�? >?P?b?t?�?�?�?�? �?�?�?OO(O:O? ^OpO�O�O�O�O�O�O �O __$_6_H_Z_l_ PO�_�_�_�_�_�_�_ o o2oDoVohozo�o �o�_�o�o�o�o
 .@Rdv��� ���o���*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4��X�j�|� ������į֯���� �0�B�T�f�J����� ����ҿ�����,� >�P�b�tφ�j�|��� ��������(�:�L� ^�p߂ߔߦ߸ߜ��� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
  �@Rdv��� ����*< N2r����� ��//&/8/J/\/ n/�/d�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�/�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�?__,_ >_P_b_t_�_�_�_�_ �_�_�_oo�O:oLo ^opo�o�o�o�o�o�o �o $6o,ol ~������� � �2�D�V�h�Lx� ����ԏ���
�� .�@�R�d�v�����~� ��П�����*�<� N�`�r���������̯ �����&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0��T�f�xߊߜ� ������������,� >�P�b�F߆���� ��������(�:�L� ^�p�����x������ �� $6HZl ~��������  2DVhz� �������/ ./@/R/d/v/�/�/�/ �/�/�/�/??�(? N?`?r?�?�?�?�?�? �?�?OO&O8OJO.? nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ `O�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�_�o�o�o, >Pbt���� ���o��(�:�L� ^�p���������ʏ܏ � ���6�H�Z�l� ~�������Ɵ؟��� � �2�D�(�h�z��� ����¯ԯ���
�� .�@�R�d�v�Z����� ��п�����*�<� N�`�rτϖ�z����� ������&�8�J�\� n߀ߒߤ߶��߬��� ���"�4�F�X�j�|� �������������� �0�B�T�f�x����� ����������, �Pbt���� ���(:L ^B������ � //$/6/H/Z/l/ ~/�/t�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�/�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O�?_*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o
_Jo\o no�o�o�o�o�o�o�o �o"4F*o<o| �������� �0�B�T�f�x�\�� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ �� ��$�6�H�Z�l� ~�������ƿؿ��� ��2�D�V�h�zό� �ϰ���������
�� .�@�$�d�v߈ߚ߬� ����������*�<� N�`�r�Vߖ����� ������&�8�J�\� n��������������� ��"4FXj| �������� 0BTfx�� �������,/ >/P/b/t/�/�/�/�/ �/�/�/??(?/8? ^?p?�?�?�?�?�?�? �? OO$O6OHOZO>? ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ pO�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�_�o�o*< N`r����� ���o�&�8�J�\� n���������ȏڏ� ���"�4�