A��*SYSTEM*   V8.2306       4/24/2014 A5  *SYSTEM*  ��AAVM_WRK_T  � $EXPOSURE  $CAMCLBDATE $PS_TRGVT   $TRGVT  $TRGHZ  $TRGDIST  $TRGW  $TRGP  $TRGR  $LENS_CENT_X  $LENS_CENT_Y  $DISTORT   $CMP_GC_P  $UTNUM  $PRE_MAST_CT   	$PRE_GRV_MST  $NEW_MAST_CT   	$NEW_GRV_MST  $STAT_RUN  $RES_ERR  $VTCP_ERR   $TRGT_ERR   $RES_ERR2  $VTCP_ERR2   $RSM_MAST_CT   	$STAT_START  $STAT_END  $STAT_ORGBK  $STAT_RSMBK  $STAT_ORGRES  $STAT_UPDT  �ABSPOS_GRP_T   $PARAM   ��ALRM_RECOV_T    $ALMRECOVENB   $ALMRECOVON   �ALMDG_T  0 $DEBUG1  $DEBUG2  $DEBUG3  $CONT_TYPE  �ALM_IF_T  D $ENABLE  $LAST_ALM d$LAST_UALM d$KALM_MAX  $LDEBUG   
 h�APCOUPLED_T  $ $APP_PROCES0  $APP_PROCES1   \�APCUREQ_T  � $SOFTPART_ID  $TOTAL_EQ  $CUR_EQNO  $PS_SPI_INDE   $SPI_INDEX  $SCREEN_NAME $APP_SIGN $APP_PROCES0  $APP_PROCES1  $TOPK_FILE 	$THKY_FILE 	$PANE_EQNO   	$DUMMY12  $DUMMY13  $DUMMY14  ��ARG_STR_T  � $TITLE $ITEM1 $ITEM2 $ITEM3 $ITEM4 $ITEM5 $ITEM6 $ITEM7 $ITEM8 $ITEM9 $ITEM10 $ITEM11 $ITEM12 $ITEM13 $ITEM14 $ITEM15 $ITEM16 $ITEM17 $ITEM18 $ITEM19 $ITEM20 �ASBN_CFG_T  8 $CNV_JNT_POS  $DATA_CMNTS  $FLAGS   $POS_CHECK  �AT_CELLSETUP 	 P $HOME_IO_PRG %$HOME_MACRO %$REPR_MACRO %$PRODRUN_SPD  $PRODRSM_SPD   �AUTOBACKUP_T 
 $ENABLE  $DEVICE $TIME   $DI_IDX  $STARTUP_BCK  $INTERVAL  $DISP_UNIT  $BCK_DO_IDX  $ERR_DO_IDX  $FR_FREE  $IN_PROGRESS  $REQ_BACKUP  $PRC_WAIT  $AUTO_BACKUP  $POFF_COUNT  $DEL_COUNT  $LOG_IDX  $DEL_TIME ? $DEL_FILE ?� $PROC_FILE ���MOTOR_COUNTE  0 $REM_COUNTS   	$REM_REV   	$BIL_REV   	��AXIS_COUNTER   $ODOMETER $NON_CMD ��AXIS_METER_T    $ODOMETER   	$NON_CMD   	��AXSCRDCFG_T  d $CARD_EXIST  $FSSB_TYPE  $CHKBD_SEL  $DIAG_REG   $SLOT_NUM  $SLOT_PREV  $DEBUG   ��BACK_EDIT_T  � $PROGRAM %$SRC_NAME %$EPT_IDX  $OPEN_ID  $DELETE_OK  $USED_TP_CRT  $BACKUP_NAME %$PS_REPLACIN   $REPLACING  $BCK_COMMENT $D_REPLACING  $SEL_PROGRAM %$DUMMY12  $DUMMY13  X�BLAL_OUT_T  , $DO_INDEX  $PS_BATALM_O   $BATALM_OR  �CFCFG_T  X $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $COMP_SWITCH  $MAX_NSETS  �CF_PARAMGP_T  � 
$WARNMESSENB  $CHKJNTLIM  $CNSTNT_CORN  $TIMEFLTRENB  $TRATIO_TB   $ACCTIME_TB1   $ACCTIME_TB2   $ORIENT_TYPE  $DEBUG  $RTSPD_SF  h�CHG_PRI_T   $TASK_ID  $PRIORITY  ��CHKPOS_T  x $CONT_FLAG  $POS_HDR  $JPOS1  $JPOS2  $JPOS3  $JPOS4  $JPOS5  $JPOS6  $JPOS7  $JPOS8  $JPOS9   	�COCFG_T  < $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $ENABLED  �CO_MORGRP_T  t $FLEN  $ANGLE  $TBA_MAG  $TBA_MAG_PRE  $TBA_MAG_MAX  $TBA_MAGAXS   	$TBA_CURAXS   	$TBA_PRVAXS   	��CO_PARAMGP_T  � $OPT_TIME  $OPT_ACC  $JACC_RRATIO  $CACC_RRATIO  $JTIME_RATIO  $CTIME_RATIO  $JVARDMAX  $CVARDMAX  $WARNMESSENB  $DEBUG  $TBA_MGN  l�CP_RSMOFST_T  @ $RO_ENABLE  $RO_MAX_ITP  $RO_NOM_DIST  $RO_NOM_SPD   ��CPCFG_T  � $GROUP_MASK  $CP_DEBUG  $CP_ENABLE  $COMP_SWITCH  $EXTRA_INT   $EXTRA_FLT   
$TF_MODE  $MD3ITPTOL  $RESUME_OFST $CP_HSTART  $T1_HSTART  $TEST   $COMP_SW2  $COMP_SW3  $COMP_SW4  ��CPDBGDEF_T  d $OUTPUT  $FILENAME )$GROUP_MASK  $DEBUGMASK  $MAXDATA  $COUNT  $TAIL  $BUFEXIST  ��CPDBG_T  � $OUTPUT  $CPIDEBUG $CPPDEBUG $MIDEBUG $MPDEBUG $MGDEBUG $MFDEBUG $SIMQSTOP  $KEEP  $PATH )$EXTRA1  $EXTRA2  L�CP_L64FIX_T  � $ENABLE  $DEC_A   $DEC_V   $DEC_CIF   $DEC_PCHO   $ADD_A   $ADD_V   $ADD_CIF   $ADD_PCHO   $DEBUG_SIM  $SIM_ADDRESS  $SIM_VAR_TYP  $SIM_AXIS  $EXTRA1  $EXTRA2  $EXTRA3  ��CP_MCRGRP_T  4 $RSM_JBF_PCT  $RSM_DEC_PCT  $RSM_OFS_PCT   �CP_MORGRP_T  � $CHNS_EMPTY  $GTF_EMPTY  $CHK_T1_SPD  $T1_FPSPD  $T1_TCPSPD  $SPEED  $T1SPDLIM  $SPEEDTOL  $JNT_VEL   	$JNT_ACC   	$JNT_JRK   	$SEGFRACTION  $RSTRT_LINE  $RSTRT_PVF  �CP_TESTDEF_T    $ENABLE_TEST  $NUM_LINES  ��CP_PARAMGP_T  D )$WARNMESSENB  $DEBUG  $ENB  $NUM_CHN  $NUM_JBFSET  $NUM_JBF  $EXT_NUM_JBF  $JBF_SIZE  $EXT_JBF_SIZ  $NUM_TF  $TF_SIZE  $EXT_TF_SIZE  $NUM_RSINFO  $JNT_VEL_LIM   	$JNT_ACC_LIM   	$JNT_JRK_LIM   	$T1SEGFL_SF  $T1GTFL_SF  $CRCMP_SWITC  $ACCLIM_SF  $JRKLIM_SF  $PSPD_SWITCH  $MAX_PSPD  $MIN_PSPD  $PSPDACC_SF  $PSPDJRK_SF  $CDCOMP_SW  $CDACC_SF  $CDJRK_SF  $CDDELTATOL  $CDDISTSF  $CDANGTOL  $CDDEVTOL  $CHKJNTLIM  $FDANG_TOL  $FDLIN_TOL  $JNTJBF_ENB  $COMP_SW  $EXTRA_INT   $EXTRA_FLT   $CP_TEST l�CP_T1_MODE_T ! � 	$ENABLE  $COMP_SWITCH  $MARGIN  $TIME_FACTOR  $SPD_LIMIT  $SLEW_RATE  $MIN_TFLEN  $EXTRA_INT   $EXTRA_FLT    \�CRCFG_T "� $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $PGDEBUG  $CR_ENHANCED  $LGORN_ENBL  $BLEND_ENB  $MAX_ARC_ANG  $RSM_RSPD_LM  $LGORN_METH  $LGORN_DBG  $LGORN_RAD  $LGORN_AZ_SP  $LGORN_ELTOL  $ROTSPDFCTR  $MAX_FP_SPD  $SMCRC_RADI  $SMCRC_RADO  $SMCRC_ARC  $ARCANGLIM  $MAXORNTCHG  $MAXSGRATIO  $CHKBMP  $RSM_TYP  $CHK_MSK  $AES_SINGTOL  �CRI_CFG_T #  $CRI_SW  �CSXC_PARAM_T $ x 	$NAME $ATTR  $NUM_CHANNEL  $IMG_HEIGHT  $IMG_WIDTH  $VT_SPACING  $DEF_ASPECT  $MIN_EXPO  $MAX_EXPO  �CUSTOMMENU_T % $ $TITLE $PROG_NAME %$OPTION  �CZ_CDCFG_T & x $ENABLE   $CD_ENABLE  $NO_HEADER  $COMP_SWITCH  $WARNMESSENB  $EXTRA_INT   $EXTRA_FLT   $CHK_SPD_SF  X�DBPXWORK_T '  $SKP_DEL    ��DBTB_CTRL_T ( � $ACRT_MODE  $MINDT_ADJ  $DELAY_CALL  $DELAY_DO  $DELAY_PLS  $RESERVED1  $RESERVED2  $RESERVED3  $NUM_IO  $DUMMY9  $DUMMY10  $�DB_DBG_T )  $DBG_PRM   
h�DPOS_DAT_T *  $X  $Y  $Z  ��LDPOS_DAT_T +  $X  $Y  $Z  \�PD_T ,  $X  $Y  $Z  L�PC_T -  $X  $Y  $Z  ��PENETRATE_T .  $X  $Y  $Z  ��DB_RECORD_T /H $CPOS *$LPOS +$DPOS_DST  $LDPOS_DST  $LINE_NUM  $ONCE_DC  $CROSS  $TASK_ID  $ENABLED_TIM  $TRIGGER_TIM  $PAUSED_TIME  $RETURNED_TI  $MMR_STATUS $CRE_NEWMON  $SIGNAL_ACT  $LAST_ACT  $PD ,$PC -$PN_AT .$PD2  $PC2  $PT  $PD_DOT_PC  $LINE_DST  $P_NUM  $GO_AWAY  $MOTION_COMP  X�DCSS_DEVICE_ 0 P $TYPE  $RBT_NUM  $SPI_IDX  $SPO_IDX  $SPI_BYTE  $SPO_BYTE  $STO  �DCSS_LS_T 1 H $STOOUT_IDX  $STOFB_IDX  $STOFB_CH  $FENCE_TYPE  $FENCE_IDX  �DCSS_PARAM_T 2 H $DOCHK_ENB  $PMCS_ENB  $LS_STOP  $LS_FENCE  $HOTSWP_TIME   t�DCSS_ELEM_T 3 T $USE  $LINK_NO  $LINK_TYPE  $UTOOL_NUM  $SHAPE  $SIZE   $DATA    ��DCSS_RBT_T 4 � $MDL_ELEM 23 
$ESTOP_DIST  $ESTOP_SPD  $CSTOP_DIST  $CSTOP_SPD  $ESTOP_JDIST   	$ESTOP_JSPD   	$CSTOP_JDIST   	$CSTOP_JSPD   	$FB_TOL   	$RBT_TYPE  $�DCS_CFG_T 5� $DISP_MENU  $LOG_ENB  $LOG_LEN  $LOG_FILE $LOG_ID  $LOG_IDMAX  $LOG_DELAY  $LOG_WRT  $LOG_INTVL  $LOG_EVENT  $TEST_PARAM1  $TEST_PARAM2  $CHK_J_TOL  $CHK_C_TOL  $SAFE_SPD  $SAFE_SPD_SV  $EXCLUDE   $SPD_ONLY   $SYS_PARAM  $PROTECT  $HI_VRC  $APPLY_WARN  $HIDE_MENU  $HI_VRC_MLT   $VRFY_ALL  $HI_MATE  $IOC_PROT  $IOC_CRC1  $IOC_CRC2  $OPI_VRC  �DCS_CRC_OUT_ 6  $START_GRP    �DCS_SGN_T 7 � 
$CURR_SIGNAT  $CURR_DATE $PREV_SIGNAT  $PREV_DATE $ANNUNC_TYP  $ANNUNC_IDX  $CUR_TIME   $LATCH_TIME   $CUR_CRC   $LATCH_CRC    d�DEFLOGIC_T 8 @ $FUNC_TITLE 	$TOTAL_NUM  $DUMMY2  $DUMMY3  $DUMMY4   �DEMO_INIT_T 9 L $DEMO_ENB  $DEMO_AU  $DEMO_DAYS  $LOAD_NUM  $DUMMY4  $DUMMY5  �EFF_AXIS_T :  $NUM  $COEFF  H�ADJ_RTRQ_T ; D $COR_TRQ   $COR_TEMP   $EFF_AXIS 2: $LIMIT  $ADJ_NUM  P�AMP_COEF_T < 0 $COEF_A   	$COEF_C  $MASK  $DUAL_MASK  �CTRL_CAB_T = @ $TRANS_A  $IDLE_PWR  $AMP_COEFB  $SV_NUM  $SV_AMP 2< �DIAG_GRP_T >8 *$VAL_SET  $TACC   	$TACC_LIM1   	$TACC_LIM2   	$RRATE_LOAD   	$VER $ANSWER  $RCC_ANS  $ADJ_RTRQ 2; $ADJ_OHTRQ   	$COPPER   	$IRON   	$BRK_PWR   	$CABLE_ACT   $CABLE_BASE   	$CABLE_LENG   	$CAB_NUM  $CTRL_CAB 2= $TRQCNS   	$TRQDWN   	$MSBAS   	$MAXTRQ   	$RRATE   	$LIFECALC   	$L10   	$N0   	$T0   	$CUR_L10   	$TCP_TYPE  $CUR_TCP $MOTN_STYLE  $FLAG  $CUR_OVC   	$CUR_HEAT   	$SUPPORT_TYP   	$ALL_SUPPORT  $CUR_TCP_X  $CUR_TCP_Y  $CUR_TCP_Z  $CUR_TCP_W  $CUR_TCP_P  $CUR_TCP_R  �DICT_CFG_T ? ` $CACHE_ENB  $CACHE_SIZE  $CURR_ONLY  $LANG_SUFFIX $LOCALE  $DUMMY5  $DUMMY6   P�DMSW_CFG_T @ 8 $KEYIMAGE  $TMS_DSB  $TMS_STAT  $TMS_INPUT    ��DOCVIEWER_T A  $DBGLVL  $CURFILE ?� 	��DPM_CFG_T B x 
$ENABLE  $DPM_INLINE  $GRP_MSK  $BEF_JBF  $DELAY  $ORI_CTL  $CUR_SCH  $MAX_SCH  $COMP_SW  $DEBUG  ��OFS_CHN_T C � $ENABLE  $OTF_DI_IDX  $CHN_TYP  $RAMP_GAIN  $SCAN_RATE  $INI_OFS  $REM_OFS  $APP_OFS  $IN_TICK  $OU_TICK  $ID  $STAT  $MAX_LIM  $MIN_LIM  $MAX_INC  $MIN_INC  $A1  $A2   4�AI_CHN_T D  $P_GAIN  $D_GAIN  $I_GAIN  $STR_CNT  $REF_CNT  $AVE_CNT  $FBK_MODE  $REF_VAL  $RAW_FBK  $CAL_FBK  $PORT_NUM  $CAL_DONE  $SLOPE  $INTERCEPT  $CUR_TICK  $LEAD_DIS  $BUF_SIZE  $BUF_CNT  $T_ADJ  $MIN_VAL  $MAX_VAL  <�BI_CHN_T E D $DI_IDX1  $DI_IDX2  $BUMP_OFS  $BUMP_RATE  $BUMP_GAIN   ��GI_CHN_T F  $DI_IDX  $SCALE   �DPM_GRP_T G � $OFS_TYPE  $OFS_FRAM  $LAST_DPM  $OFS_ACCU  $OFS_ABS  $OFS_CARRY  $CTL_RATE  $INT_LINE  $OFS_LINE  $DAT_RDY  $OFS_STAT  $SND_TYPE  $TRK_MODE  $SYNC_DI  $OFS 2C 	$AI_CH 2D 	$BI_CH 2E 	$GI_CH 2F 	H�DPM_SCH_T H 0 $GRP_MSK  $COMMENT $DPM_ON  $GRP 2G ��DPM_IN_T I 8 $LINE_NUM  $DELAY  $OFS_X  $OFS_Y  $OFS_Z  ��DRC_CFG_T J D $HOST1 !$HOST2 !$HOST3 !$HOST4 !$HOST5 !$EMAIL_ENABL  <�DSBL_FAULT_T K  $ENABLE  $MAX_COUNT  8�DTREC_T L, $DTREC_ENB  $SAMPLE_ITP  $BUF_SIZE  $FILE_SIZE  $DEVICE_NAM $SUBBUF_SIZ  $SPC_FILE  $DTREC_ON  $DTSAV_ON  $FILE_ACCESS  $PC_ACCESS  $SYSTIME   P$DTSAV_ENB  $ORDER  $DSB_BUFSIZ  $ENB_BUFSIZ  $OTTASK_MOD  $DP_ALM_ID  $DP_ALM_GRP  $DP_ALM_AXS  $DEF_MAXBUF  x�DYN_BRK_T M 0 $DI_IDX  $DO_IDX  $BRK_MSK  $FLTR_IF  (�ENC_STAT_T N� $ENC_COUNT  $ENC_ROS_TIK  $ENC_RATE  $ENC_AVERAGE  $ENC_ENABLE  $ENC_DSPSTAT  $ENC_SPCSTAT  $ENC_SIM_ON  $ENC_SIM_SPD  $ENC_VALUE  $ENC_HEAD  $ENC_MULTIPL  $ENC_STOPPED   $ENC_THRESH  $ENC_EXISTS  $ENC_HSDI  $ENC_ABSCNT  $INCTRAVDIST  $INCTRAVCNTS  $INCTRAV_DO  $CONVSPD_GO  $INCTRAVRES  $ENC_BUFFER   d$ENC_ATR_AXS  $SC_GRP_NUM  $ENC_COMERCT  $ENC_FBCMPCT  �ENETMODE_T O 8 $FULL_DUPLEX  $SPEED  $ACD_ENABLE  $THROTTLE  ��ER_NOAUTO_T P D $NOAUTO_ENB  $NOAUTO_NUM  $PS_NOAUTO_C   $NOAUTO_CODE    8�ER_NOALM_T QH *$NOALMENBLE  $NOALM_NUM  $ER_CODE1  $ER_CODE2  $ER_CODE3  $ER_CODE4  $ER_CODE5  $ER_CODE6  $ER_CODE7  $ER_CODE8  $ER_CODE9  $ER_CODE10  $ER_CODE11  $ER_CODE12  $ER_CODE13  $ER_CODE14  $ER_CODE15  $ER_CODE16  $ER_CODE17  $ER_CODE18  $ER_CODE19  $ER_CODE20  $ER_CODE21  $ER_CODE22  $ER_CODE23  $ER_CODE24  $ER_CODE25  $ER_CODE26  $ER_CODE27  $ER_CODE28  $ER_CODE29  $ER_CODE30  $ER_CODE31  $ER_CODE32  $ER_CODE33  $ER_CODE34  $ER_CODE35  $ER_CODE36  $ER_CODE37  $ER_CODE38  $ER_CODE39  $ER_CODE40  ���ER_OUTPUT_T R � $OUT_NUM  $IN_NUM  $PLCWARN  $GRP_STR  $ERROR_NUM  $FAC_NUM  $SEV_NUM  $PARM1_NUM  $PARM2_NUM  $DUMMY9  $DUMMY10  $DUMMY11   ��EXT_SET_T S < $ENABLE  $DI_TYPE  $DI_NUM  $DO_TYPE  $DO_NUM  8�FDR_GRP_T TT $VEL_MOD   	$VEL_CNT   	$REM_LIFE2   	$OVM_RATE   	$OVA_RATE   	$TROV_RATE   	$DTAV_RATE   	$DTMX_RATE   	$DTMIN_RATE   	$MOT_RATE   	$DIAG_INDX_R   
$DIAG_INDX_I   $DG_MAXT   	$DG_T0   	$RATED_TRQ   	$DRIVE_TYPE   	$GEAR_RATIO2   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$Z_MCMD   	��FEATURE_T U , $NAM ? $MOD ? $VER ? $MEC ?   �FILECOMP_T V  $TPP  $VARIABLE  `�FILE_SETUP2_ W 4 $FILE_TDC_SC  $FILE_TV_SEC  $FILE_TVC_SC   X�FILE_BACK_T X T $FILE_NAME )$PROG_NAME %$FUNC_CODE  $MODIFIER  $COMMENT %$FUNC_PTR    ��FMR2_GRP_T Y $VEL_ROT  $VEL_LIN  $VEL_MOD   	$K_LIFE   	$NTR_LIFE   	$EFF_RATE   	$ROT_INRT   	$TROV_MAX   	$T_LIFE_0  $RATED_TRQ   	$LIMIT_FUNC  $ACC_LMT   	$DRIVE_TYPE   	$GEAR_RATIO2   	$DGCLFR   	$DGDYFR   	$DGLDEC   	$DG5T0   	$DG_MAXT   	$DG_T0   	$�FMR_CFG_T Z  $TROV_MAX   T�FSSB_CFG_T [ P $FSSB_LINE   $EX_FSSBLINE   $FSSB1_AXES  $FSSB3_AXES  $FSSB5_AXES  �GRAVC_GRP_T \ � 
$MODE_SW  $SPCONS   	$DEBUG1  $DEBUG2   	$GRV_STATUS  $BKUP_NO116   	$POFF_NO116   	$GRVCMP_SW  $GRVMST_LOOP  $MST_SMT_LEN   ��MOTYPE_E ]       �TERMTYPE_E ^      �ORIENT_E _    �ޠ�SM_PROFILE_E `    �b8�TA_PROFILE_E a       �UPR_T b� -$MOTYPE ]$TERMTYPE ^$SEGTERMTYPE ^$DECELTOL  $USE_CONFIG  $USE_TURNS  $ORIENT_TYPE _$UFRAME $UTOOL $SPEED  $ROTSPEED  $CONTAXISVEL  $CNSTNT_PATH  $CNSTNTPTHJT  $SEG_TIME  $USE_CARTACC  $USEMAXACCEL  $USERELACCEL  $USETIMESHFT   $USE_PATHACC  $USE_SHORTMO  $SM_PROFILE  `$TA_PROFILE  a$ACCEL_OVRD  $TIME_SHIFT  $ACCU_NUM   $PAYLOAD  $DYN_I_COMP  $PATHRES_ENB  $RESERVE1   $CNT_SHORTMO  $EXT_SPEED  $CNT_ACCEL1  $CNT_ACCEL2  $CRCCOMPENB  $ASYMFLTRENB  $USE_WJTURNS  $EXT_INDEP  $CARTFLTRENB  $CNT_SPEEDUP  $CNT_DYN_ACC  $MAX_SPEED  $USERELPSPD  $PSPD_OVRD  $ORNT_MROT  0�GRSMT_GRP_T c  $GRV_SW  $GRV_PARAM   ��HOST_CFG_T d � $COMMENT $PROTOCOL 	$PORT $OPER  $STATE  $MODE $REMOTE $REPERRS  $TIMEOUT  $PATH e$STRT_PATH e$STRT_REMOTE $USERNAME e$PWRD_TIMOUT  $SERVER_PORT  $USE_VIS_PRT  ��HOSTENT_T e 4 $H_NAME !$H_ADDRTYPE  $H_LENGTH  $H_ADDR !�ERR_MASK_T f H $SSC_MASK1  $SSC_MASK2  $SSC_MASK3  $SSC_MASK4  $SEV_MASK  4�HSCD_MNG_T g $COLL_MODE  $THRESHOLD  $DO_ERR  $DO_ENABLE  $MACRO_REG  $STND_CD  $AUTO_RESET  $UPD_GROUPS  $PARAM_VERID 	$PARAM119   	$PARAM120   	$PARAM121   	$PARAM122   	$PARAM123   	$PARAM124   	$PARAM125   	$ACT_RATIO  $SAVED119   	$SAVED120   	�HSCD_GRP_T h $ $COL_DET_OFF  $HSCD_PRM_ID  $�HTTP_AUTH_T i ( $OBJECT !$NAME $TYPE  $LEVEL  �HTTP_T j � $ENABLE  $ENAB_DIAGTP  $ENAB_SPART  $DBGLVL  $KRL_TIMOUT  $HITCOUNT  $BG_COLOR $ENAB_TEMPL  $TEMPLATE $COMMENT $RSS_INUM  �HWR_CONFIG_T k H $MAINCPU  $VISIONCPU  $SPARE1  $SPARE2  $SPARE3  $SPARE4  h�IBGN_CFG_T l $CMP_WAIT  $MAX_PNUM1  $MAX_PNUM2  $FWD_TOL_LOC  $FWD_TOL_ORT  $FWD_TOL_EXT  $FWD_TOL_ANG  $BWD_TOL_LOC  $BWD_TOL_ORT  $BWD_TOL_EXT  $BWD_TOL_ANG  $BWD_RTN_SPD  $UF_DATA  $DBG_MASK  $TEMP_MGN  $LIN_N_CNST  $END_TOL_LOC  $STATUS  $RECDAT_SEND    �IBGN_ERRIO_T m @ $REC_IO_TYP  $REC_IO_NUM  $EXE_IO_TYP  $EXE_IO_NUM   0�IBGN_EXEC_T n ( $SCHEDULE   $FILE_P   $BWD_FLG     H�IBGN_FIL_T o @ $EXE_MD  $EXE_OPN  $EXE_BACK  $REC_TRANS  $REC_ACC  ��IBGN_FTP_T px $FTP_CTAG  $AUTO_TRANS  $IGNR_COMER  $FTP_STAG  $SM_STAG  $SM_CTAG  $SM_SPORT  $SM_CPORT  $N_PCSOFT 	$N_RECFL1 	$N_RECFL2 	$N_RECFL3 	$N_EXEFIL $N_FLEXT1 $N_CONDFL 	$N_FLEXT2 $N_SPTXT1 $N_SPTXT2 	$SEQ_VAR  $SNS_NUM  $SNS_CNST  $FOLDER $RECS_PRG %$RECS_TMO  $RECE_PRG %$RECE_TMO  $SM_DBG  $AUTO_START  $RESERVE  \�IOLNK_T q 8 $RACK  $SLOT  $INPUT_N  $OUTPUT_N  $OPTION  ��IOSLAVE_T r  $INPUT_N  $OUTPUT_N   ��IO_DEF_ASG_T s T $LOG_TYPE  $LOG_NO  $NUM_PORTS  $RACK  $SLOT  $PHY_TYPE  $PHY_NO    ��IO_UOP_CFG_T t ` $UOP_TYPE  $IN_RACK  $IN_SLOT  $IN_STRTPT  $OUT_RACK  $OUT_SLOT  $OUT_STRTPT   x�UJR_GRP_T u � $FINE_OVRD  $JOGFRAME $FINE_DIST  $J7_GROUP  $J8_GROUP  $J7_AXIS  $J8_AXIS  $J7_LABEL $J8_LABEL $J7_GRAPHIC Q$J8_GRAPHIC Q$DSB_J7J8  $DSBL_KEY   �KAREL_CFG_T v 0 $CONV_ENABLE  $CONV_CTRL  $CONV_FLAGS  	��LGCFG_T w � $ENABLE  $OUT_SW  $LG_SIZE  $EV_SIZE  $MR_SIZE  $SG_SIZE  $FD_SIZE  $MI_SIZE  $ER_SIZE  $MP_SIZE  $MG_SIZE  $PE_SIZE  $LG_MODE  $EV_MODE  $MR_MODE  $SG_MODE  $FD_MODE  $PE_MODE  $EX_RSCH_FIL $COMP_SW  L�LN_DISP_T x ` $HIDE_LINE_N  $DISP_MENU  $HIDE_PARLN  $HIDE_DAULN  $HEAD_PARENT $HEAD_DAUGHT   ��LOGBOOK_T yt B$NUM_ER_ITM  $NUM_ER_TYP  $NUM_REC_TYP  $NUM_SCRN_FL  $NUM_DIO  $SRAM_MARGIN  $DRAM_MARGIN  $OPTION  $LOG_ER  $LOG_ENT  $LOG_SEL  $LOG_WIN  $LOG_MENU  $LOG_JGMU  $LOG_MNCHG  $LOG_FNKEY  $LOG_JGKY  $LOG_PRGKEY  $LOG_UFKY  $LOG_OVRKY  $LOG_FWDKY  $LOG_HLDKY  $LOG_STPKY  $LOG_PRVKY  $LOG_ENTKY  $LOG_ITMKY  $LOG_RSTKY  $LOG_HELPKY  $LOG_OVR  $LOG_CRD  $LOG_STEP  $LOG_GRP  $LOG_SGRP  $LOG_UF  $LOG_UT  $LOG_FILE  $LOG_WTRLS  $LOG_PGCHG  $LOG_SETPOS  $LOG_TPKY  $LOG_DIO  $LOG_STMD  $LOG_FOCUS  $LOG_PRGEXE  $LOG_TUIKEY  $IMG_ENT  $IMG_SEL  $IMG_WIN  $IMG_FNKY  $SAVE_FILE 	$SCRN_FL  $SCRN_NO_ENT  $ANALOG_TOL  $AVAILABLE  $CLEAR_ENB  $DCS_HI1  $DCS_HI2  $DCS_HO1  $DCS_HO2  $DCS_SI  $DCS_SO1  $DCS_SO2  $DCS_OPTION  $IGNR_SAVE  $FNKEY_FLTR  $DCS_DEV  �LOG_BUFF_T z 0 $TITLE $SIZE  $MEM_TYPE  $VISIBLE   �LOG_STAT_T { 0 $TICK  $SPD  $POS1  $POS2  $POS3   �LOG_DCS_T | � $ENABLE  $SPD_TOL  $OUTPUT_TYP  $OUTPUT_IDX  $GRP_NUM  $POS_TYP  $AXIS_NUM  $STOP_READY  $STOP {$ESTOP {$CSTOP {$ESTOP_DIFF {$CSTOP_DIFF { �LOG_DIO_T } L $RACK  $SLOT  $MOD_TYPE  $PORT_TYPE  $START_PORT  $END_PORT  �LOG_SCRN_FL_ ~  $SP_ID  $SCRN_ID   �MCSP_T  � $CLDPOP_ENB  $TRQLIM_ENB  $JOGLIM_ENB  $CLDPOP_FLG  $CLDGRP_FLG  $CLDREL_FLG  $CLR_CLDFLG  $JOGLIM_FLG  $ORGJOG_OVR  $COMP_SW  $RESERVE1  $RESERVE2  $RESERVE3  H�MCSP_GRP_T � � 	$JOGLIM_OVR  $TRQLIM_FLG  $SV_PTLIM   	$ORG_PTLIM   	$ORG_RCLMC   	$RESERVE1  $RESERVE2  $RESERVE3   	$RESERVE4   	 �MISC_GRP_T � d $HPD_TRQ   	$DSTB_MAX   	$DSTB_MIN   	$DSTB_MAXENB   	$DSTB_MINENB   	$DSTB_EXCESS  $e��MISC_MSTR_T �  $HPD_ENB  ���MISC_SCD_T � H $DSTB_MAX_A   	$DSTB_MIN_A   	$DSTB_MAXENB   	$DSTB_MINENB   	��MKCFG_T � \ $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $MO_CONFLICT  $MO_REQUIRED  $DEBUG  L�MLTARM_CFG_T �  $NUM_ARMS  $GROUP   U�MLT_GRP_DO_T � � $TP_ENABLE  $JOG_GROUP  $LOCKED_ARM  $CRNT_TYPE  $CRNT_INDX  $PRG_ROUT_P  $JOG_ROUT_P  $PRG_DO_TYPE   $PRG_DO_INDX   $JOG_DO_TYPE   $JOG_DO_INDX    �MNDSP_MST_T � ` $DISP_ENABLE  $DISP_EDCMD  $DISP_INAUTO  $DISP_RSMDIS  $DISP_IS_ON  $MODE_GRP   *P�MNDSPPSTL_T � 4 $LOCTOL  $ORIENTTOL  $EXTTOL  $ANGTOL   		��MODAQ_CFG_T � d $ON_LINE  $MF_FLAG  $MI_FLAG  $GRP_NUM  $STARTLOG  $ENDLOG  $LN_MASK  $SUPPORT   ��FX_TRIGGER_T � � 	$START_MODEL  $START_STEP  $START_PROG %$STOP_MODEL  $STOP_STEP  $STOP_PROG %$AXES  $DATA_TYPE  $DATETIME  ��MODEM_INF_T � t $MDM_INIT )$MDM_INIT1 )$MDM_RESET )$MDM_HANGUP )$MDM_DIAL )$MDM_ANSWER )$MDM_STATUS )$MDM_IDENT )��MOR_GRP_SV_T �  $CUR_SV_ANG   	�ARMLOAD_T �  $ARMLOAD   X�ARMLOAD_P_T �  $ARMLOAD_P    ��MRR2_GRP_T �� $ARM_PARAM   d$CALIB_MODE  $GEAR_PARAM   2$SPRING_PAM   <$RLIBSW01  $RLIBSW02  $ABC_FLAG  $MD_J2SECT   $MD_J3SECT   
$MD_J1SPCONS   P$MD_J2SPCONS   P$MD_J3SPCONS   P$MD_CUR_K   $MD_CUR_J2  $MD_CUR_J3  $SV_OFF_TIM2   	$CSKPLIM_ENB  $CSKPLIM_LIN  $CSKPLIM_JNT   	$QSKPLIM_ENB  $QSKPLIM_LIN  $QSKPLIM_JNT   	$EXT_AZIM   $EXT_ELEV   $SERVOCMPTOL   	$ARMLOAD 1� $ARMLOAD_X 1� $ARMLOAD_Y 1� $ARMLOAD_Z 1� ��INTERACT_T �  $INTERACTION   	��INTRAC_N_T �  $INTRAC_NUM   	��INTRAC_D_T �  $INTRAC_DIV   	��DH_EXTRA_T � 0 $VALID  $X  $Y  $Z  $W  $P  $R  |�MRR_GRP_T �H �$BELT_ENABLE  $CART_ACCEL1  $CART_ACCEL2  $CIRC_RATE  $CONTAXISNUM  $PS_EXP_ENBL   $EXP_ENBL  $JOINT_RATE  $LINEAR_RATE  $PATH_ACCEL1  $PATH_ACCEL2  $PATH_ACCEL3   $PROCESS_SPD  $PROC_SPDLIM  $CNT_ACC_MGN  $DDACC_RATIO  $FWP_TIME1  $FWP_TIME2  $ACCEL_RATIO  $DECEL_RATIO  $PPABN_ENBL  $ROTSPEEDLIM  $SPEEDLIM  $SPEEDLIMJNT  $DEF_MAXACCE   $USE_CAL  $SPIN_CTRL  $SYN_ERR_LIM   $SYNC_GAIN   $SYNC_OFFSET   $MOUNT_ANGLE  $COLLINEAR  $COINCIDENT  $ACCEL_TIME1   	$ACCEL_TIME2   	$ENCSCALES   	$EXP_ACCEL   	$PS_INPOS_TI   $INPOS_TIME   	$JNTVELLIM   	$JNT23_UPLIM  $JNT23_LOWLI  $LOWERLIMS   	$LOWERLIMSDF   	$MASTER_POS   	$MIN_ACCTIME   	$MOSIGN   	$MOT_SPD_LIM   	$PERCH    	$MOVERRLIM    	$PERCHTOL    	$STOPERLIM   	$STOPTOL   	$SERVO_CTRL  $PS_SV_OFF_A   $SV_OFF_ALL  $SV_OFF_ENB   	$SV_OFF_TIME   	$UPPERLIMS   	$UPPERLIMSDF   	$TRKERRLIM  $PAYLOAD  $PS_MAX_PAYL   $MAX_PAYLOAD  $AXISINERTIA   	$AXISMOMENT   	$MAX_AMP_CUR   	$ACCEL_PARAM   $MAX_PTH_ACC  $MRRDUM2   $PS_BCKLSH_C   $BCKLSH_COUN   	$MOVER_GAIN   	$MOVER_SCALE   	$MOVER_OFFST   	$CLALM_TIME  $TSMOD_TIME  $CHKLIMTYP  $SNGLRTY_STP  $INPOS_TYPE  $JOG_TIME_M  $MIN_ACC_UMA  $MIN_ACC_UCA  $ACC_SCL_UCA  $SLMT_J1_LW   $SLMT_J1_UP   $SLMT_E1_LW   $SLMT_E1_UP   $SLMT_J1_NUM  $SLMT_E1_NUM  $PS_SPCCOUNT   $SPCCOUNTTOL   	$SPCMOVETOL   	$SHORTMO_MGN  $MIN_ACC_CMC  $EXTACCRATIO  $CN_GEAR_N1  $CN_GEAR_N2  $SFLT_ERLIM   	$SV_CTRL_TYP   	$PS_CARTMO_M   $CARTMO_MGN  $MIN_CAT_UMA  $MIN_ACC_SHM  $GEAR_RATIO   	$EXP_JOG_ACC   	$PS_ARMLOAD   $ARMLOAD   $ACC_PA_UMA  $ACC_PC_UMA  $AXIS_IM_SCL  $PS_MOT_LIM_   $MOT_LIM_STP  $JG_FLTR_SCL  $JOGACCRATIO   $TORQUE_CONS   	$MIN_PAYLOAD  $DECOUP_MGN   $DECP_MGN_WR   	$PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $FFG_MGN_J2  $FFG_MGN_J3  $DVC_AC0_MAX   	$DVC_AC1_MAX   	$DVC_ACC_MAX   	$DVC_ACC_MIN   	$DVC_JRK_MAX   	$DVC_JRK_MIN   	$SV_DBL_SMT  $SV_MCMD_DLY  $SV_GRV_X  $SV_GRV_Y  $SV_GRV_Z  $SV_DH_D   	$SV_DH_A   	$SV_DH_COSA   	$SV_DH_SINA   	$SV_LNK_M   	$SV_LNK_X   	$SV_LNK_Y   	$SV_LNK_Z   	$SV_LNK_IX   	$SV_LNK_IY   	$SV_LNK_IZ   	$SV_Z_SIGN   	$SV_DMY_LNK   	$SV_DH_COSTH   	$SV_DH_SINTH   	$SV_THET0   	$LNK23Z  $LNK23X  $LNKCBZ  $LNKCBX  $CB_MASS  $CB_IX  $CB_IY  $CB_IZ  $LNKSBY  $LNKSBX  $LNGTSB  $SPCNS  $ARMLOAD_X   $ARMLOAD_Y   $ARMLOAD_Z   $DUTY_ENB   	$DUTY_PARAM1   	$DUTY_PARAM2   	$QSTOP_TOL   	$NE_ENB  $LINK_TYPE   	$ARMLOAD_NUM   	$DH_THETA0   	$DH_THETA   	$DH_D   	$DH_A   	$DH_ALPHA   	$LINK_M   	$LINK_SX   	$LINK_SY   	$LINK_SZ   	$LINK_IX   	$LINK_IY   	$LINK_IZ   	$DH_VD   	$DH_VA   	$DH_VALPHA   	$LINK_VM   	$LINK_VSX   	$LINK_VSY   	$LINK_VSZ   	$LINK_VIX   	$LINK_VIY   	$LINK_VIZ   	$DH_HD   	$DH_HA   	$DH_HALPHA   	$LINK_HM   	$LINK_HSX   	$LINK_HSY   	$LINK_HSZ   	$LINK_HIX   	$LINK_HIY   	$LINK_HIZ   	$DH_OTHETA   	$DH_OD   	$DH_OA   	$DH_OALPHA   	$LINK_OM   	$LINK_OSX   	$LINK_OSY   	$LINK_OSZ   	$LINK_OIX   	$LINK_OIY   	$LINK_OIZ   	$FLINK_BX   	$FLINK_BY   	$FLINK_BETA   	$SPBALANCE_K   	$SPLENGTH_0   	$SPACT_X   	$SPACT_Y   	$SPACT_Z   	$SPFULC_X   	$SPFULC_Y   	$SPFULC_Z   	$INTERACTION 1� 	$AUTO_SNGSTP  $T1T2_SNGSTP  $CART_2ND_TI  $JNT_2ND_TIM   	$LC_QSTP_ENB  $CP_CUTOFFOV  $CP_MINSEG  $MASTREV_ENB  $MASPOS_DIFF   	$INTRAC_NUM 1� 	$INTRAC_DIV 1� 	$OBS_DIST  $SV_PARAM   2$MIJNTCHKLMT  $LCHWARN_ENB  $ABC_PARAM   $MECH_MASK  $MECH_TYPE  $AXS_MAP_NUM  $AXS_MAP   	$DH_EXTRA 1� 
$AXS_COUPLE   	$PS_ROBOT_CR   $ROBOT_CRC   ��MSK_CE_GRP_T � P $T1_USERCART  $T1_USERJNT   	$T1_CARTVEL  $T1_JNTVEL   	$T1_WARNING  �MTCOM_CFG_T �  $CNC_NO  $NORES_TIMEO  �OPWORK_T �, $SYSBUSY  $SOPBUSYMSK  $TPBUSYMSK  $UOPBUSYMSK  $INTPRUNNING  $INTPPAUSED  $INTPMASK  $OPT_OUT  $UOP_DISABLE  $OUTIMAGE   $OP_PREV_IMG   $OP_INV_MASK   $ORGOVRDVAL  $USER_OUTPUT   $PS_ENBL_ON   $ENBL_ON  $MLT_RBT_ENB  $PMC_EDT_MSK   $NOALM_MSK  $DUMMY19  ��OVRDSLCT_T � x $OVSL_ENB  $SDI_INDEX1  $SDI_INDEX2  $OFF_OFF_OVR  $OFF_ON_OVRD  $ON_OFF_OVRD  $ON_ON_OVRD  $DUMMY  �$�OVRD_SETUP_T � @ $OVRD_NUM  $OVERRIDE   
$OVRD_NUM_S  $OVERRIDE_S   
 �TRACECTL_T � H $TASK_STATUS  $TRC_TOP_IDX  $TRC_BTM_IDX  $TASK_ID  $DUMMY4  �TRACEDT_T � D $EPT_INDEX  $LINE_NUM  $FILE_OFST  $EXEC_TYPE  $LINE_ST  �TRACEUP_T � @ $TRC_UPDATE  $DISP_PXNN  $DUMMY2  $DUMMY3  $DUMMY4  ��PG_CFG_T � $SUBTASKNUM  $NUM_TASKS  $JMPWAIT_UPR  $JMPWAIT_LOW  $FAST_MODE  $RCVFAIL_CNT  $WAITREL_CFG  $ACC_CTRL  $CNT_CTRL  $IGNR_PLS  $DBTB_STPTYP  $BWD_CFG  $RESUME_CFG  $IGPAUS_PRI  $MTNLN_CFG  $PAUS_RTN  $RESERVE1  $RESERVE2  ��PG_DEFSPD_T � L $AP_DEF_SPD  $AP_DEF_UNIT  $DUMMY4  $APSP_PREXE  $DLY_LASTPS   ��PING_T � 0 $TIMEOUT  $DATALEN  $NPACKETS  $DEBUG  �PIPE_CFG_T � h $ARSIZE   $FILEDATA   $SECTORS  $FORMATTER  $RECORDSIZE  $MEMTYPE  $FORMAT  $AUXWORD   ��PLID_CFG_T �  $COMP_SWITCH   H�MAX_PLD_CAL_ � $ $AA  $BB  $CC  $DD  $EE  �CALC_RESULT_ � � $PAYLOAD  $PLD_J3ARM  $INERTIA4  $INERTIA5  $INERTIA6  $MOMENT4  $MOMENT5  $MOMENT6  $COMB_LOAD4  $COMB_LOAD5  $COMB_LOAD6  $PUB_INRT4  $PUB_INRT5  $PUB_INRT6   #��PLID_GRP_T �P H$PI_ENB  $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $ARMLOAD3  $ROB_TYPE  $DATA_NUM  $SPEED_HIGH  $SPEED_LOW  $DEFSPD_HIGH  $DEFSPD_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DEFACC_HIGH  $DEFACC_LOW  $SAMPLE_TIME  $SAMPLE_HIGH  $SAMPLE_LOW  $MOV_AXIS   	$MOV_POS1   	$MOV_POS2   	$MOV_DEF1   	$MOV_DEF2   	$ROT_INERTIA   	$MAX_VEL_HI   	$MIN_VEL_HI   	$MAX_ACC_HI   	$MIN_ACC_HI   	$MAX_VEL_LOW   	$MIN_VEL_LOW   	$MAX_ACC_LOW   	$MIN_ACC_LOW   	$GAMMA   	$STOP_DATA  $GETDATA_FIN  $ID_RESULT   
$CALIBRATE  $PI_DEBUG  $HIDAT_V_MAX   	$HIDAT_V_MEA   	$HIDAT_A_MAX   	$HIDAT_A_MEA   	$LWDAT_V_MAX   	$LWDAT_V_MEA   	$LWDAT_A_MAX   	$LWDAT_A_MEA   	$CALC_TYPE  $MTN_CALCTYP  $CHKER_VER $PDCK_RB_TYP  $I_FACTOR   $MAX_PAYLOAD  $MAX_INERTIA   $MAX_MOMENT   $COMB_LOAD   $MAX_PLD_CAL �$IM_SRCH_DT  $WARN_DISP  $WARN_LEVEL  $OVER_LEVEL  $CALC_RESULT �$PAMSWFLG  $AMLD_SCRN  $DUMMY69  $DUMMY70  $DUMMY71    �PLID_SV_T �P $CUR_SCRN  $CUR_GROUP  $PS_SAVE_DON   $SAVE_DONE  $NO_RECOVER  $RESULT_SAV   
$PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  $ARMLOAD1  $ARMLOAD2  $DO_DEFAULT  $MOV_POS1   	$MOV_POS2   	$SPEED_HIGH  $SPEED_LOW  $ACCEL_HIGH  $ACCEL_LOW  $DO_DEF_POS   x�PLIM_GRP_T � � $MAX_PYLD  $AXISINERTIA   	$AXISMOMENT   	$AXIS_IM_SCL  $PS_LIM_WT_S   $LIM_WT_SCL  $LIM_INR_SCL   $LIM_MNT_SCL   $LIM_CL_SCL   $PLD_MODE  $DUMMY10  $DUMMY11  ��PLMR_GRP_T � � $PYLD_ENB  $WMR_ENB  $ANGLE  $PLMR_AA  $PLMR_BB  $PLMR_CC  $PLMR_DD  $PLST_ANG   
$COMP_SW  $MAX_XY_LOC  $MAX_Z_LOC  �PLST_GRP_T � p $COMMENT $PAYLOAD  $PAYLOAD_X  $PAYLOAD_Y  $PAYLOAD_Z  $PAYLOAD_IX  $PAYLOAD_IY  $PAYLOAD_IZ  �PL_RES_G_T � | $PAYLOAD  $SAVMOMENT4  $SAVMOMENT5  $SAVMOMENT6  $SAVINERTIA4  $SAVINERTIA5  $SAVINERTIA6  $EST_RESULT   ��PL_RES_V_T �  $PL_RES_G_P   �PMON_QUE_T � 8 $QCOUNT  $QTHRESHOLD  $QHYSTERESIS  $QUEUE_UP  �PM_GRP_T � � $ACC_TIME1  $ACC_TIME2  $POS_ERR_LIM  $ROT_ERR_LIM  $ENABLED  $DBG_MASK  $COMP_SWITCH  $BWD_ACC1  $BWD_ACC2  $JVEL_RATIO  $REWIND_NUM  $GTF_ACC1  $GTF_ACC2  �POCFG_T �   $PODEBUG  $OVERRUN_TOL   ��PODATA_T � P $OVERRUN_CNT  $CUR_INDEX  $PROGRAM_ID   2$LINE_NO   2$OVERRUN_ITP   2�POINFO_T �  $CUR_INDEX  $INFO   ��POIO_T � ( $SLEQ_NUM  $IO_TYPE  $IO_INDEX  ��POS_EDIT_T � � 	$LOCK_POSNUM  $HIDE_MENU  $HIDE_POSNUM  $AUTO_RENUM  $COPY_POSDAT  $AUTO_RENUM2  $RMV_MANRENM  $COPY_POSTYP  $CPRUT_ENB   �PRGADJ_T � h $X_LIMIT  $Y_LIMIT  $Z_LIMIT  $W_LIMIT  $P_LIMIT  $R_LIMIT  $SPEED_ADJ  $NEXT_CYCLE  ,�PRGNS_CFG_T � � $ALGO_VER  $NYQ_FREQ  $WIN_TYPE  $WIN_SIZE  $OVERLAP  $FREQ_LIM  $MIN_NUM  $CREATED  $VERIFY  $PROGNAME %$CREATE_GP  $STATUS_GP  $DEBUG  $MAILTIME  $MAILEVENT  $LASTMAIL  �PRGNS_ELEM_T � � $ENABLE  $FEASIBLE  $AXIS  $PS_ELEM_NUM   $ELEM_NUM  $ROT_RATIO  $MAX_FREQ  $THRE_REL  $THRE_ABS  $DEGRAD_LVL  $DEGRAD_BASE  $DEGRAD_RATE  $UPD_DATE $BASE_DATE ��PRGNS_GRP_T � X $ELEM 2� $MIN_ANG   	$MAX_ANG   	$BASE_ANG   	$LAST_MOD   	$BASE_MOD   	 "��PRGNS_PREF_T � ( $GRIDLINES  $BARS_NUM  $STYLE  ,�PROTOENT_T �  $P_NAME !$P_PROTO  �PROXY_CFG_T � � $LIST_PORT  $PROXY_ENB  $PROXY_SRV )$PROXY_PORT  $DIRECT_1 )$DIRECT_2 )$DIRECT_3 )$DIRECT_4 )$DIRECT_5 )$DIRECT_6 )$DIRECT_7 )$DIRECT_8 )��PF_DATA_T �   $VALUE  $GROUP  $AXIS  0�PF_CFG_T �| $ENABLE  $PROG_NAME %$CUR_GROUP  $RAN_GROUPS  $START_TYPE  $TOTAL_TIME  $TOTAL_PWR  $INS_PWR  $REGEN_PWR  $INS_REGEN  $EXE_DATE $DATA_TYPE  $RES_NAME %$MONTR_RATE  $D_PWR_SUP  $D_PWR_REG  $RV_LIM1  $RV_LIM2  $DEGREE  $REFRESH  $OVERRIDE  $RV_HRS_DAY  $RV_DAYS_YR  $MAXSIZE  $SUMMARY 2� $CONFIG_SET  $SUPPORT  $LAST_RUN  ��PF_PREF_T � 4 $GRIDLINES  $BARS_NUM  $DATA_TYPE  $STYLE  �PSSAVE_T � $MC_FOLDER 	$SLAVE_SAVE  $START_MULTI  $SLAVE_LOAD   $LOAD_DEV  $KEEP_HNADDR !$KEEP_HRADDR !$KEEP_CCOMM $KEEP_CPROT 	$PS_KEEP_COP   $KEEP_COPER  $KEEP_CSTATE  $KEEP_CREMOT $KEEP_CTIMEO  $KEEP_CSREMO $KEEP_CUNAME e$KEEP_CHPWD  $KEEP_SBMSK !<�PSSAVE_GRP_T � , $FLANGE  $SYNC_FLANGE  $SYNC_MST_CN  �PS_CONFIG_T � � $DB_IMMTRIG  $DA_IMMTRIG  $DB_NOTRIG  $DA_NOTRIG  $TCLAMP_WARN  $USE_DYNSPD  $MAX_SEARCH  $NUM_PSMOTN  $DB_MARGIN  $RESOLUTION  $COMP_MASK  $PX_STARTED  $SCAN_READY  $SCAN_ALIVE  �PS_CP_CFG_T �  $ENB  $REF_MODE  ��PS_CP_GRP_T � � 
$ENB  $REF_MODE  $FLANG_VALID  $FLANG_TICK  $FLANG_TRANS $PREVI_TRANS $UTOOL_VALID  $UTOOL_TRANS $FKSOL_FP  $SEG_COUNTER  ��PS_ITEM_T � � $BASE_DIST  $TUNE_MSEC  $MN_LEN  $ITEM_LINE  $ITEM_DONE  $TRIGGERED  $STOP_TRIG  $NG_ITEM  $CLAMPED  $PARAM1  $PARAM2  $PARAM3  $ML_ACT_P  $MN_CODE   �PS_MOTION_T ��  $OWNER_TID  $G0  $PS_DONE  $PG_STATUS  $DB_STATUS  $DA_STATUS  $DB_MIN_DIST  $DA_MAX_DIST  $PARENT_NAME %$CHILD_NAME %$PARENT_LINE  $SCAN_COUNT  $SEG_STARTED  $SEG_COUNTER  $SCAN_ABORT  $PARENT_EPT  $CHILD_EPT  $PRV_VALID  $PRV_DB_DIST  $PRV_DA_DIST  $PRV_VEC   $PRV_TICK  $BASE_SPEED  $DEST_VALID  $DEST_VEC   $UT_TRANS $MMR_P  $MODONE  $NEXT_MODONE  $SMH_MASK  $NUM_ITEM  $ITEM 2� h�PWRUP_DLY_T �   $DELAY_TIME  $SY_READY   8�QSKIP_GRP_T � � $ERROR_CNT2   	$QSKP_ERRCNT   	$QSKP_CURANG  $QSKP_CURAN1  $QSKP_CURAN2  $QSKP_CURAN3  $QSKP_CURAN4  $QSKP_CURAN5  $QSKP_CURAN6  $QSKP_CURAN7  $QSKP_CURAN8  $QSKP_CURAN9  �J2RED_T � 4 $EXD_RTQ  $EXD_ITP  $EXD_PRG  $EXD_LINE  ��RDCR_GRP_T � � $RMAX_TORQUE   	$RMIN_TORQUE   	$THRES_TORQ   	$RGEAR_RATIO   	$WARN_FLG   $COMP_SW  $RESERVE   	$SPC_ITP  $NUM_EXD  $J2TH2ND  $J2RED 1� ��REFPOS11_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS21_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS31_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS41_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS51_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS61_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPOS71_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  `�REFPOS81_T � l $COMMENT $ENABLED  $ATPERCH  $DOUT_TYPE  $DOUT_INDX  $PERCHPOS   	$PERCHTOL   	$HOMEPOS  ��REFPSMSK_T �  $MAXREFPOSEN    ���REMOTE_CFG_T � 4 $REMOTE_TYPE  $REMOTEIOTYP  $REMOTEIOIDX   ��REPOWER_T �  $FLAG  ��RESTART_T � , $FLAG  $DSB_SIGNAL  $STARTUP_CND   ��RS232_CFG_T � � $COMMENT $DEVICEUSE  $SPEED  $PARITY  $STOPBITS  $FLOWCONTROL  $TIMEOUT  $CUSTOM  $AUXTASK  $INTERFACE  $STATUS  '��RSCH_T � @ $OLD_SPEC_SW  $FREEFROMSIZ  $TARGET_DIR 	$UPDT_MAP   �RSPACE_T �� !$COMMENT $USAGE  $ENABLED  $IN_EXTERIOR  $ENTRY  $ENT_SIGN_ON  $PRIORITY  $PRIORWRK  $DOUT_TYPE  $DOUT_INDX  $DIN_TYPE  $DIN_INDX  $FRIEND_GRP  $UFRAM_NUM  $UTOOL_NUM  $MYHOLD  $LENGTH_VTEX  $FIRST_VTEX   $SECND_VTEX   $UFINV_POST $MARGIN  $WAITING  $FIRST_VTX2   $SECND_VTX2   $G2ENTRY  $G1ENT_INTR  $G2ENT_INTR  $PRE_UFRAM  $NO_USE_DI  $HOLD_REQ  $CSPACE_NUM  $CUR_TCP   $PRE_TCP   ��GP_STATUS_T � @ $IN_USE  $SPACE_NUM  $PRIORITY  $STATUS1  $STATUS2  ��COM_SPACE_T �X $USE_MLT_CTN  $H_PRIORITY  $IN_CONTROL  $IN_SPACE_GP  $WT_SPACE_GP  $USE_GP  $DEADLOCK_GP  $DELAY_CNT1  $DELAY_CNT2  $GP_STATUS 2� $DOUT1_TYPE  $DOUT1_INDX  $DOUT2_TYPE  $DOUT2_INDX  $DOUT3_TYPE  $DOUT3_INDX  $DIN1_TYPE  $DIN1_INDX  $DIN2_TYPE  $DIN2_INDX  $EXT1  $EXT2  $V1   $V2   $V3   �GP_HOLD_T � � $STATUS  $GP_MSK  $SPACE_NUM  $CSPACE_NUM  $REQ_GRP  $PS_RATE   $RATE   $INT_POS   $ACT_POS   $PRD_POS   $S1  $S2  $S3  $S4   �RSPACEG_T � 0 $COM_SPACE 2� $GP_HOLD 2� $SPARE_INT   
 �RSPACESR_T � � $SR_ENB_TYP   $RUNNER_AXS  $HAND_LNGTH  $HAND_THICK  $FLIP_ENB  $INTFERENCE  $HAND_IF_CHK  $HANDI_TYPE  $HANDI_INDX  $SR_G1POS   $SR_G1POS_IN   $SR_G1ANG   $SR_G1ANG_JF   $SR_PRM   	�RTCFG_T � � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $RSM_RTCP  $INLINE_WRST   $TBC_PTH_CMP  $DRTCP_ENB  $LDR_SP_RATE  $LDR_RSP_RAT  $COMP_SWITCH   
�RV_DATA_T �  $DATETIME    	$VALUE    	�RV_DATA_GRP_ �  $DATA  2� �SCR_T �	| �$ITP_TIME  $NUM_GROUP  $NUM_TOT_AXS  $NUM_DSP_AXS  $JOGLIM  $FINE_PCNT  $COND_TIME  $MAXNUMTASK  $KEPT_MIRLIM  $MAXPREMTN  $MAXPREAPL  $PRE_EXE_ENB  $NUM_SYS_MIR  $NUM_PG_MIR  $BRKHOLD_ENB  $ENC_AXIS    $ENC_TYPE    $NUM_GP_MADE  $NUM_RLIBSOC  $NUM_MOTNSOC  $DUMMY158  $SV_CODE_OPT  $SFSPD_OVRD   $COLDOVRD  $COORDOVRD  $TPENBLEOVRD  $FENCEOVRD  $JOGOVLIM  $SFJOGOVLIM  $RUNOVLIM  $SFRUNOVLIM  $MAXNUMUFRAM  $MAXNUMUTOOL  $LCHDLY_TIME  $RECOV_OVRD  $JOGWST_MODE  $JOGLIMROT  $MOTN_PC_RUN   @$RESETINVERT  $OFSTINCVAL  $FWDENBLOVRD  $TPMOTNENABL  $PREV_CTRL  $MAX_PRE_FDO  $PRE_MB_CMP  $MB_DSBL_MSK  $MB_DSB_MSK2  $SVSTAT  $UPDATE_TIME  $JG_DSBL_MSK  $NUM_PG_AMR  $MB_LD_MSK  $MOTN_LD_MSK  $MOTN_LD_MK2  $AMP_TYPE   T$CAP_AMP_DIS   T$HBK_MAP_ENB  $HBK_IO_TYPE  $HBK_IO_IDX  $PPA_MAP_ENB  $PPA_IO_TYPE  $PPA_IO_IDX  $MOTN_LD_IDX   @$DVC_DBG  $DVC_ENB  $DVC_MODE  $DVC_MODE1  $DVC_MODE2  $DVC_MODE3  $DVC_C_RATIO  $INTASK_OVRU  $DSP_TYPE  $CABINET_TYP  $NE_MODE  $PG_DSBL_MSK  $JOG_AUX_ENB  $SUBCPU  $NE_SIN_RESO  $UPDATE_MAP1  $UPDATE_MAP2  $UPDATE_FLAG   $HW_C1_TIME1  $HW_C1_TIME2  $ATR   �$UNITTYPE   �$ATRATTRIB   �$NE_CYCLE  $NECA_OVRUN  $FLTR_2_FIX  $STARTUP_CND  $DSB_SIGNAL  $LPCOND_TIME  $CHK_CH_SCTM  $F_ATR   �$F_UNITTYPE   �$F_ATRATTRIB   �$FSSB_STAT   �$CHAIN_TIME  $CHAIN_STAT  $CHAIN_RSDN  $DSP_MAP_ENB  $IDX_TBL_MSK  $PROC_CTRL  $TEMPER_LIMS   T$FSSB1   $FSSB2   $FSSBDIAGENB  $RAILACC_ENB  $SMCR_LOADED  $DUMMY159  $PS_DSP_TYPE   $DSP_TYPE2  $PRC_DSP   $PRC_CD_ID 	$MOTN_FUNC   $INTRINS_TP  $DIAG_FUNC  $TRANS_NUM   T$TRANS_MAX   T$TRANS_WARN   T$CBLCUR_MAX   T$CBLCUR_A   T$CBLCUR_B   T$CBLCUR_WARN   T$DAC_TRANS   T$DAC_CBLCUR   T$CLDET_PT  $CLDET_AXS   $PS_CLDET_TI   $CLDET_TIME   $CE_RIA_SW  $SAFE_SPD  $SAFE_ROTSPD  $T2_LOCK_ENB  $DSB_MOINIT  $MAX_DF_LEN  $MPDT_TIMLMT  $FAST_HRDYON  $ORG_PTH_RSM  $DAC_LMT  $MULSELENB  $UPDATE_MAP3   $JCOLDOVRD  $JTPENBOVRD  $JFENCEOVRD  $FAN_ALMLVL  $FAN_WRNLVL  $HARDTYP_MAP  $COMP_SW   2$SHADOWRECS  $SHADOWTIME  $FANSTOP_TIM  $BRK_ECO_ENB  $AUTATR_STAT  $AUTO_SBRIDX  $AUTO_DSPIDX  $AUTO_ATRIDX   $AUTO_AMPINF   �$AUTO_AMPCUR   �$REGTYPE  �AX_OFS_T �  $X  $Y  $Z  0�SCR_GRP_T �� �$NUM_SEG   $NUM_PT   $ARM_TYPE  $DUMMY121  $ARM_TYPE_B  $NUM_AXES  $NUM_ROB_AXS  $NUM_RED_AXS  $WRST_AXIS_S  $WRST_AXIS_E  $SYNC_M_AXIS  $SYNC_S_AXIS  $WRIST_TYPE  $HW_STRT_AXS  $AXISORDER   	$DUMMY122  $BRK_NUMBER   	$DUMMY123  $DD_MOTOR   	$ROTARY_AXS   	$LOADRATIO   	$CONFIG_MASK  $LINK_LENGTH   $EXT_ORDER   $DUMMY124  $EXT_XYZ_MAP   $DUMMY125  $EXT_OFFSET   $EXT_LENGTH   $ROBOT_ID $ROBOT_MODEL 	$ROBOT_FILE 	$ROBOT_INT  $SV_CODE_ID $JOGLIM_JNT   	$COORD_MASK  $OP_BRK_NUM   	$DUMMY126  $USE_TBJNT  $USE_TBCART  $NUM_DUAL  $DUMMY127  $PS_TURN_AXI   $TURN_AXIS   $AXS_AMP_NUM   	$FLEXTOOLTYP  $AXS_XYZ_MAP   	$DUMMY128  $OFST 1� 	$KINEM_ENB  $DUMMY129  $PS_UPDATE_M   $UPDATE_MAP  $TORQCTRL  $DSP_NUM   	$DUMMY130  $PS_M_POS_EN   $M_POS_ENB  $M_DST_ENB  $MOVE_DST  $MCH_POS_X  $MCH_POS_Y  $MCH_POS_Z  $MCH_POS_W  $MCH_POS_P  $MCH_POS_R  $MCH_ANG   	$MCH_SPD  $DST_MIR_P  $DPOS_DST  $DST_POS_X  $DST_POS_Y  $DST_POS_Z  $DSP_ERCNT   	$PS_DEST_DAT   $DEST_DATA_P   $ROBOT_FUNC  $PROC_AXS   	$DAC_MODE  $DAC_AXMODE   	$DAC_RATE1   	$DAC_RATE2   	$DAC_RATE3   	$DAC_RATE4   	$DAC_RATE5   	$DAC_RATE6   	$DAC_RATE7   	$DAC_RATE8   	$DAC_RATE9   	$DAC_RATE10   	$DAC_LMT1   	$DAC_LMT2   	$DAC_LMT3   	$DAC_LMT4   	$DAC_LMT5   	$DAC_LMT6   	$DAC_LMT7   	$DAC_LMT8   	$DAC_LMT9   	$DAC_LMT10   	$DAC_DEBUG   $FUNC_SW   $FUNC_VAL   $ABC_ENB  $HBK_ENBL  $MV_DIAG   
$ABC_MODE1  $ABC_MODE2  $ABC_MODE3  $ABC_MODE4  $ABC_MODE5  $ABC_MODE6  $ABC_MODE7  $ABC_MODE8  $ABC_MODE9  $SAFE_JNTSPD   	$ROBOT_LABEL $DSP_NUM_FLG  $GROUP_NUM  $COMP_SW   $AMB_TEMP  $DSP_STRT_AX  $TOT_SBR_NUM  $TOT_DSP_NUM  $TOT_ATR_NUM  $TANDEM_SUB   	$DSP_ORDER   	$ATR_ORDER    $AMPINF_ORDR    $AMPCUR_ORDR    $FIX_ORNT_WR  �SERVENT_T � $ $S_NAME !$S_PORT  $S_PROTO !��SERV_MRA_T � d $DATETIME  $ERR_CODE  $SAFETY_ST  $IMP_VEL   	$IMP_TOQ   	$ANGLES   	$DIST_TOQ   	 T�SERV_REC_GRP � p $TOTAL  $BIN_V1T1   	$BIN_V1T2   	$BIN_V2T1   	$BIN_V2T2   	$MRA_REC 1� 
$MRA_IDX  $WCA_REC 1� 
��SERV_RV_T �  $OVER_LIMIT   	 �SERV_OCCUR_T �  $ERR_CODE  $COUNTER  ��SHELL_CFG_T � 5$JOB_BASE  $RSR_ENABLE   $NUM_RSR   $RSR1_NAME %$RSR2_NAME %$RSR3_NAME %$RSR4_NAME %$RSR5_NAME %$RSR6_NAME %$RSR7_NAME %$RSR8_NAME %$JOB_ROOT %$CONT_ONLY  $USE_ABORT  $RSR_ACKENBL  $INVERT_CHK  $UOP_SEL_STA  $RSR_ACK_PUL  $COM_TIMEOUT  $PNS_ENABLE  $SHELL_NAME %$START_MODE  $TPFWD_KAREL  $ERR_REPORT  $OPTIONS  $QUE_ENABLE  $PRODSTARTYP  $CSTOPI_ALL  $SHELL_EXT  $SEL_TYPE  $EXT_SEM1  $EXT_SEM2  $MAINT_STYL  $ISOL_ENB  $DI_CHKTRIG  $PROD_MODE  $INIT_TMO  $MANRQ_TMO  $EXTEND_ENB  $KEYSWITCH  $STARTCHKTYP  $HEARTBEATMS  $PERM_LEVEL  $TEMP_LEVEL  $USTART_FT  $START_SIG  $DO_HOME_SOP  $REFPS_PR_ID  $DIS_STRTCHK  $CUSTOM  $E_RECOV_MSK  $SET_IOCMNT  $CSTOPI_ALL2   l�SHELL_CHK_T � D $ENABLE  $RESUME  $PROMPT  $ERRPOST  $FORCE  $WARN   T�SHELL_COMM_T � @ $FUNC  $STATUS  $PARM1  $PARM2  $PARM3  $PARM4   p�SMB_HDDN_T �  $BLOB    �SNPX_ASG_T � 0 $ADDRESS  $SIZE  $VAR_NAME %$MULTIPLY  �SNPX_PARAM_T � � $TIMEOUT  $SNP_ID 	$NUM_ASG  $NUM_CIMP  $NUM_FRIF  $VERSION  $STATUS  $DISP_INFO  $MODBUS_ADR  $NUM_MODBUS  $MODBUS_PORT   ��SSR_T � x $SINGLESTEP  $DUMMY7  $SGLSTEPTASK   &$STEPTASKNUM  $STEPSTMTTYP  $STPSEGTYPE  $BWDSTEP  $SHOWSTMTTYP  �SVDT_GRP_T �� �$DATA00   	$DATA01   	$DATA02   	$DATA03   	$DATA04   	$DATA05   	$DATA06   	$DATA07   	$DATA08   	$DATA09   	$DATA0A   	$DATA0B   	$DATA0C   	$DATA0D   	$DATA0E   	$DATA0F   	$DATA10   	$DATA11   	$DATA12   	$DATA13   	$DATA14   	$DATA15   	$DATA16   	$DATA17   	$DATA18   	$DATA19   	$DATA1A   	$DATA1B   	$DATA1C   	$DATA1D   	$DATA1E   	$DATA1F   	$DATA20   	$DATA21   	$DATA22   	$DATA23   	$DATA24   	$DATA25   	$DATA26   	$DATA27   	$DATA28   	$DATA29   	$DATA2A   	$DATA2B   	$DATA2C   	$DATA2D   	$DATA2E   	$DATA2F   	$DATA30   	$DATA31   	$DATA32   	$DATA33   	$DATA34   	$DATA35   	$DATA36   	$DATA37   	$DATA38   	$DATA39   	$DATA3A   	$DATA3B   	$DATA3C   	$DATA3D   	$DATA3E   	$DATA3F   	$DATA40   	$DATA41   	$DATA42   	$DATA43   	$DATA44   	$DATA45   	$DATA46   	$DATA47   	$DATA48   	$DATA49   	$DATA4A   	$DATA4B   	$DATA4C   	$DATA4D   	$DATA4E   	$DATA4F   	$DATA50   	$DATA51   	$DATA52   	$DATA53   	$DATA54   	$DATA55   	$DATA56   	$DATA57   	$DATA58   	$DATA59   	$DATA5A   	$DATA5B   	$DATA5C   	$DATA5D   	$DATA5E   	$DATA5F   	$DATA60   	$DATA61   	$DATA62   	$DATA63   	$DATA64   	$DATA65   	$DATA66   	$DATA67   	$DATA68   	$DATA69   	$DATA6A   	$DATA6B   	$DATA6C   	$DATA6D   	$DATA6E   	$DATA6F   	$DATA70   	$DATA71   	$DATA72   	$DATA73   	$DATA74   	$DATA75   	$DATA76   	$DATA77   	$DATA78   	$DATA79   	$DATA7A   	$DATA7B   	$DATA7C   	$DATA7D   	$DATA7E   	$DATA7F   	 +��SVPRM_UPD_T �  $PRM   
��SVGUN_CT_T � ` $OUTPUT_ENB  $INPUT_ENB  $GROUP_NUM  $AXIS_NUM  $GO_VALUE  $GI_VALUE  $IO_SCALE  �SYSLOG_T � � $SIZE  $MODE  $STATUS  $ADDRESS  $DATA_SIZE  $COMP_VALUE  $STOP_MODE  $CURR_VALUE  $FLOG_ID_LO  $FLOG_ID_HI  $FLOG_ID_IN  $FILE_OUT  $FILE_NAME $ID  p�SYSLOG_SAV_T � h $SAVE_BLCKS  $SAVE_TASKS  $SAVE_D_CPU  $SAVE_D_SIZ  $SAVE_D_ADD  $FILE_OUT  $FILE_NAME x�SYSTEM_TIMER � p 
PWR_TOT  PWR_LAP  SRV_TOT  SRV_LAP  RUN_FLG  RUN_TOT  RUN_LAP  WIT_FLG  WIT_TOT  WIT_LAP  ��TBC_ACC_T �X -$ACC_LEN1  $ACC_LEN2  $ACCEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT   	$M_STAT  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $AC_ACC  $JK_ACC  $VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AAL1  $AAL2  $AAL3  $AAL4  $AAL5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM   <�TBCCFG_T � ` $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $TBC_STAT   $TC 2� $TBC_DEBUG  �TBCSG_GRP_T � \ $ENABLE  $APPRC_SCL   
$OPEN_SCL   
$CLOSE_SCL   
$CLS_MINF2   
$CLS_MINACC   
�$$CLASS  ������       �$$VERSION  ������  ���$AAVM_WRK 2 ������ 0  �5�                                �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            @  �                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            _POS�                                                 	 	                                     ���� 	                                     ����                                                       	                                                               �5�                            HZ �                                                 	 	                                     ���� 	                                     ����                                                       	                                                             �$ABSPOS_GRP 1������� <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �$ACC_MAXLMT        ��   ��$ACC_MINLMT        ��    �$ACC_PRE_EXE        ��    �$AC_UPDATE  �����������$ALARMRECOV ������   �        �$ALMDG ������                �$ALM_IF ������    d                                                                                                       d                                                                                                         , 
                                         �$ANGTOL  ������� 	 A   A   A   A   A   A   A   A   A   �$APPLICATION ?������� 
 HandlingTool          
V8.20P/A2             
88150                 
3367298              
1829               �0
V8.20P/A2          �  7DE3/A2               	80604.015             FRL                  H2                   ��$AP_ACTIVE      ����   �$AP_AUTOMODE         �    �$AP_CHGAPONL         �   �$AP_COUPLED 1�������                                                                  �$AP_CUREQ 1������   T                                          	           	            	 ���                                          	           	            	 ���       �Handling      HT           	           	HTTHKY     	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ���                                          	           	            	 ����$AP_CURTOOL      ����   �$AP_DO_CLEAN         �    �$AP_DO_CLENM  �������                                                                                                                          �$AP_DSPDRYRN         �    �$AP_HIDE  ������� @                                                                                                                                                                                                                                                                 �$AP_MAXAPP         �   �$AP_MAXAX          �    �$AP_PLUGGED      ����   �$AP_PRC_DSBM  �������                                  �$AP_PROC_DSB         �    �$AP_SEGF_CHK         �    �$AP_SEG_CHKM  �������                                                                                                                          �$AP_SELAP  ������� @                                                                                                                                                                                                                                                                �$AP_TOTALAX      ����    �$AP_USENUM  �������   �$ARG_STRING 1������� 
�MENUS             
MENU_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                I/O SIGNALS       Tryout Mode       Input Simulated   Output Simulated  OVERRIDE = 100    In cycle          Prog Aborted      Tryout Status     	Heartbeat         MH Fault          MH Alert            n                  n                  n                  n                  n                  n                  n                  n                  n                  n                TOOL              
TOOL_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                WORK              
WORK_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                POS               	POS_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                DEV               	DEV_ITEM1           n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PALT              
PALT_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                GRIP              
GRIP_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                USER              
USER_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                PREG              
PREG_ITEM1          n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                  n                �$ARG_WORD ?	�������  	$         	[         	]         	�          	�          �$ASBN_CONFIG �������           �$ASCII_SAVE            �    �$ATCELLSETUP 	�������%  OME_IO                               %MOV_HOME                              %MOV_REPR                                      �$AUTOBACKUP 
�������    FRA:\                                             '`                       �                 15/12/03 07:06:06         �                          �                          �                          �                            ��                                                                                                                                       ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      ��                                                                                                                                      �  RA:\_BACKUP_\ATBCKCTL.TMP DATE.DT                                                                                                �$AUTOINIT         �    �$AUTOMESSAGE        �   �$AUTOMODE_DO         �   �$AUTOMODE_OV         �   �$AUTOPAUSPOS !��������  (7��ɓ]>��������M��W��V�            )�B��3                                9�B�r�                                I�                                    (O����������������������������(O����������������������������(O����������������������������(O�����������������������������$AUTOPPOSTSK  �������                              �$AUTOUPDTMOD         d�   �$AXIS_COUNT 1������   �  � 	 �+} �6 n-y��� K����w             	  1j? c�T J�q ,�� 8�W BcR             	                                      	 J������� �'L_�|�             	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXIS_METER 1������   �  P 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$AXSCRDCFG 1������  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �$BACKGROUND         �   �$BACKUP_NAME 	�������	BACKUP    �$BACK_EDIT 1������� 
 �%-BCKEDT-                              %UP021                                 �     ��%-BACKUP-                              �    �                        %-BCKEDT-                              ��%-BCKED2-                              %  AKRO050                              �       %-BACKU2-                                    �                        %  BCKED2-                              ��%-BCKED3-                              %                                       ���      %-BACKU3-                                    �                        %-BCKED3-                              ��%-BCKED4-                              %�                                      ���      %-BACKU4-                                    �                        %-BCKED4-                              ��%-BCKED5-                              %�                                      ���      %-BACKU5-                                    �                        %-BCKED5-                              ��%-BCKED6-                              %�                                      ���      %-BACKU6-                                    �                        %-BCKED6-                              ��%-BCKED7-                              %�                                      ���      %-BACKU7-                                    �                        %-BCKED7-                              ��%-BCKED8-                              %                                       ���      %-BACKU8-                                    �                        %-BCKED8-                              ��%-BCKED9-                              %                                       ���      %-BACKU9-                                    �                        %-BCKED9-                              ��%-BCKCRT-                              %�                                      ���      %-BACCRT-                                    �                        %-BCKCRT-                              ���$BCK_NO_DEL         �   �$BGE_UNUSEND         �   �$BLAL_OUT �������  �   �$BWD_ABORT         �    �$BWD_ITR_RTN         ��   �$BWD_NONSTOP         �   �$CE_OPTION         �   �$CE_RIA_ID         �   �$CFCFG �������                      �$CF_PARAMGP 1�������                                                                                                     C�  C�  C�  C�  C�  D  D  D  D  D  D  D   D%  D*  D/  D4  D9  D>  DC  DH    D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D�� D��         ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�                                                                                                      C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�    C|  C�  C�  C�� C�� C�� C�� C�� C�  C�  C�  C�  C�  Cʀ CЀ Cր C܀ C� C�  C�          ?�  �$CHECKCONFIG         �    �$CHG_PRI 1�������         ��������������������������������������������������������������������������������������������������������������������$CHKPAUSPOS 1�������  ,    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    ������������������������������    �������������������������������$COCFG �������              �$CO_MORGRP 2�������  �   ^B�0�?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  �$CO_PARAMGRP 2�������  ,       ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�         ?   ?   ?�  ?�     K   K       ?�  �$CPCFG ������          a�m                                                                                   
                                            ����                @                                 �`        �$CPDBG ������        )cpmidbg                                      �   �  :�  +�  +�       )cpmpdbg                                      �     �  J  K       )midbg                                        �     �   �   �       )mpdbg                                        �     �   -   .       )mgdbg                                        �     �  g  h       )mfdbg                                     ���������                    )ud1:                                              �$CPDBGDEF ������       )ud1:cpdbgbuf.txt                             �                    �$CP_L64FIX ������                                                                                                                                                                                                                                                                                                                                                                                                                                               �$CP_MCRGRP 2������     d   d   d   d   d   d   d   d   d   d   d   d�$CP_MORGRP 2������  �                 ?��;CH  BH   	 B��'B�S�B�E�B�LB�ECD�             	 C~�C�kC�.VC�S�Cˇ�D2a"             	 EI�EQEc/rE���Eis�E�|~            ?�     7                         CH  BH   	 F8�R                                 	 Ip=�                                 	 Mh.                                ?�     7                         CH  BH   	 FYQO                                 	 I�{�                                 	 M88�                                ?�     7                         CH  BH   	                                      	                                      	                                     ?�     7    �$CP_PARAMGRP 2 ������ <                        b  �     b  x    	 C  C� C� C�  C4  DH               	 D&��Da  DS3FZfĎ�F*tf             	 D�0 E �fD���GB� E�p GA��            ?�  >�33 ;��@   @�         n   @   @�   5�@�  @   ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    ������                    ~      d  �      d  x    	 E�                                   	 H��                                  	 J;�                                 ?�  >�33 ;��?�  @          n   @   @�     	@   @�  ?�  ?@  A�  ?       =L��<#�
                                                    �������$CP_RSMOFST ������                  �$CP_T1_MODE !������     G   
?@      ;��
                                               �$CP_TESTDEF ������           �$CRCFG "�������                             C4  A�             �   x   A�  Cz  B�  CH  B�  CH  C  @�     -       :d�
�$CRI_CFG #�������   �$CRT_DEFPROG %�������%�                                      �$CRT_INUSER         �    �$CRT_KEY_TBL  ������   	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������͓�����������������������������耇���������������������$CRT_LCKUSER         �    �$CRT_USESTAT         �    �$CR_AUTO_DO        ��    �$CR_INDT_ENB         �   �$CR_T1_DO        ��    �$CR_T2_DO        ��    �$CSTOP         �   �$CSXC_PARAM 2$������ 
 8
SONY XC-56                    �  �@���?�     ( АSONY XC-HR50                  �  �@���?�     ( АSONY XC-HR57                  �  �Aff?�     ( А�                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �                                                      �$CTRL_DELETE         �   �$CT_POPUP             �    �$CT_QUICKMEN         �    �$CT_SCREEN �������kcsc  �$CT_USERSCRN �������c_sc  �$CUSTOMMENU 1%������  <               %                                                          %                                       ���               %                                       ����              %�                                      ����              %�                                      ���Start SM Comm %IBSCMANS                              ���End SM Comm   %IBSCMANE                              ���User Cancel   %UCANCACT                              ���
User Reset    %URESACT                               ����              %�                                      ����              %�                                      ����              %�                                      ���Zange         %ZG_MENUE                              ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���VAG_KONFIG.   %VW_MENUE                              ����              %�                                      ���VAG-Dateien   %DATEIEN                               ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���
Macro Step tt %MSK_STAT                              ���Wait Monitor  %SHTPEST                               ����              %�                                      ����              %�                                      ���CYCLE POWER   %PWDCYCLE                              ���
POWER DOWN    %	PWD_MAINT                             ����$CUST_MANUAL         �   �$CZCDCFG &�������            	                                              ?|(��$DBCONDTRIG         �   �$DBLOVRD_ENB         �   �$DBNUMLIM        d�   
�$DBPXWORK 1'�������                                                                                                                          �$DBTB_CTRL (�������                ���$DB_AWAYTRIG      GCP �=��
�$DB_AWAY_ALM         �    �$DB_CONDTYP         �   �$DB_DBG 1)�������  , 
               ,  	     �  *        
                                        �$DB_MINDIST      GCP �@�  �$DB_MONTIME        ��  ��$DB_MONTYP         
�   �$DB_MOTNEND         �   �$DB_RECORD 1/�������  �                        G�O�G�O�   .            U��U��    U��EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   /            U��U�+    U�EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�               U�U�=    U�7EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�               U�7U��          XECUTING

 ����                                                                  G�O�                                    G�O�G�O�               Uc�UgK    Ug_EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   (            U6cU8�    U7EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   ,            U7�U9�    U8%EXECUTING

 ����                                                                  G�O�                                    G�O�G�O�   0                              TOPPING
�O&n�                                                                  G�O�                                    G�O�G�O�                                  XECUTING
�S��� 1                                                                G�O�                                    G�O�G�O�                                  CANCELLED
    - l                                                                G�O�                                    G�O�G�O�                                                190                                                                G�O�                                    G�O�G�O�                                                201                                                                G�O�                                    G�O�G�O�                                                )
$                                                                G�O�            �$DB_TOLERENC      B�  �=L���$DCSS_DEVICE 10������                                                                                                                                                                                                                            �$DCSS_LS 11������                                                                                                                                                                  �$DCSS_PARAM 2������                 �$DCSS_RBT 24������ 8 
 <                  D	�       ��  �                                    B�                D�         ��                   Cπ       B�  C      �A� C                        C\        C�  �H                                    C        B   �H      İ@ �H                        CH            �           �   �          c                                                     c                                                     c                                                     c                                              C���Dz  D	;Dz   	 BG��A{�A���@ͤ�AIXA�Z�             	 B�  B�  B�  B�  B�  CH               	 B[��A�  A�C�A陚A�  B>ff             	 B�  B�  B�  B�  B�  CH               	  �R O|O ��� P   P   P                   
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                          
 <       c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                     c                                                               	                                      	                                      	                                      	                                      	                                         �$DCS_CFG 5�������          dMC:\DCSL%04d.CSV                     c                   �    A   A   CH  Cz                                                                                �            �   �   �   �   �   �   �            �`iMU��    �$DCS_CRC_OUT 6�������                  �$DCS_C_FSI ?������ �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_FSO ?������ P �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$DCS_C_RPI ?������  �                      �                      �                      �                      �$DCS_C_RPO ?������  �                      �                      �                      �                      �$DCS_SGN 7�������e+u�12-JUN-24 17:06   ���03-DEZ-15 07:06            IK(�IK(�H<=H<=                    e+u��,s��i�ZX�_                  �$DCS_VERSION �������V3.3.2            �$DEFLOGIC 18�������  	�          ���	�          ����	�          �����$DEFPROG_ENB         �   �$DEFPULSE         ��   �$DEF_ACCLIM        ��   ��$DEF_WRSTJNT         �����$DEMO_ENB            �    �$DEMO_INIT 9���������������� ���$DEMO_OPT_SL ?	������   � 
 	R575      	R745      	R746      	R747      	R750      	R751      	R752      	�          	�          	�          �$DEMO_OPT_TO  ������   � 
                                         �$DEV_INDEX         d�   �$DEV_PATH A�������A\KJLTVL111120R01\ 01\  \ \ 20\ JE\ OLGE123_SEPARADO\              �$DHCP_CLNTID ?�������  �                  �                  �$DIAG_GRP 2>������ �   
 	 F?h FR� FR� Eu  Eu  D�               	 B�  B�  B�  B�  B�  B�               	 B�  B�  B�  B�  B�  B�               	 CVV�Cc� C���CH�kCAUSB�"�            f362 678901234567890          �  BG�B�Bz�B�B
Q�B��BA���A��A�
=                  @�  A   Ap  A�  A�  A�  B  B   B4                        ������       
  B'33B#�BB�B��B�BBz�B
=Bz����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  B!�B=qB�RB�Bp�B�B��B�
B�RA������������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A�(�A���A��A�Q�A��HA~�RAw�Ap  AhQ�A`Q����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A�
=A�(�A���A�\)A��
A�=qA}�Aup�Amp�AeG����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
  A��HA��
A��RA��A�=qA��HAz�HAs�
Al��Ae����������      @�  A   Ap  A�  A�  A�  B  B   B4  ���������  ������������       
 	 B
Q�B��Bp�A��HA��
A�=q             	 =}�=m�h=m�h>8Q�>8Q�>8Q�             	 7��8b08b07�Ŭ7�Ŭ7�Ŭ             	 @ʏ\@ʏ\@ʏ\@�p�@�p�@�p�              @�  Ah  A�       	 <#�
<#�
<49X=#�
=#�
=#�
             	 ;#�
;#�
;#�
;��
;��
;��
                 �>���C�  <(�U     4 	 @�  @�  @�  @���@���@���            A@     ?     	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	 ?+�?G+?G+?#�
?#�
?#�
             	 ��G���G���G���G���G���G�             	 B�  B���B���B   B   B                	 B�  B�  B�  A�  A�  A�               	 CVW
Cc� C��
CH�)CAT{B�#�             	                                	   p  p  p  p  p  p             	 Ap  Ap  Ap  Ap  Ap  Ap               	 E�  E�p E�p D�  D�  DD               	                                         8�>�C?�'�5~�����5i�]��>��|�4���x�,D���D���   0        	                                      	                                      	                                  �x�,D���D���´  B4�Bp      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                      	                                      	                                      	                                      	                                     12345678901234567890          �                                                                                                                      ������          ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������  ���������������������������������������  ���������������������������������������  ������������������ 	                                      	                                      	                                      	                                                        	                                      	                                           �                  4 	                                                  	 ������������������������������������ 	 ������������������������������������������������  4 	 ������������������������������������ 	 ������������������������������������ 	 ������������������������������������ 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                         8�                                                             	                                      	                                      	                                                                 �$DICT_CONFIG ?�������          eg      ���$DISTBF_TTS         
�   �$DISTBF_VER        
�   �$DMAURST         �    �$DMSW_CFG @������               �$DOCVIEWER A������     	 ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  �$DPM_CFG B������                          
        �$DPM_SCH 2H������ 
�   Schedule 1            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 2            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 3            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 4            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 5            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 6            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 7            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 8            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 9            �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz     Schedule 10           �                     ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz                       ?�                               	 H          ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?             ?�  ?�                              A       >L��    ?   ?    	 TA   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz  A   A   A      
   
   
                      ?�                             Dz   	         =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A           =L��?�  A    	     Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz      Dz  �$DPM_SIM 2I������                                                                                                                                                          �$DRC_CFG J�������!�                                  !�                                  !�                                  !�                                  !�                                     �$DSBL_FAULT K�������        �$DSBL_GPMSK         ��    �$DTDIAG L������            UD1: 678901234567890                         P                                                                                                                                                                                                                                                                                                                                              �               @   �$DTRECP L������            
UD1:                                          P                                                                                                                                                                                                                                                                                                                                              �               @   �$DUMP_OPTION  �������    �$DUTR_CFG      ����   �$DUTR_CPMES      ����   �$DUTY_TEMP  È�3B�  �A�  �$DUTY_UNIT         �    �$DYN_BRK M�������        �$ED_SIZE    '   �  x �$ED_STATE         �    �$EMGDI_STAT      ���     �$ENC_STAT 1N������  �                                                                     
                 d                                                                                                                                                                                                                                                                                                                                                                                                                                 ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ������������������������������������������������������������������ d ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        �$ENETMODE 1O�������                                            �$ERROR_PROG %�������%�                                      �$ERROR_TABLE  �������  �������������������������������������������������������������$ERRSEV_NUM       ��   �$ER_AUTO_ENB         �    �$ER_NOAUTO P�������          *�  *�  *�  *�  *�  +                                                        �$ER_NOHIS         �    �$ER_NO_ALM 1Q�������  �         *�  *�  *�  *�  +                                                                                                                                            �$ER_OUT_PUT 2R�������    @�                ����$ER_SEV_NOAU  �������                 �$ETCP_VER !�������!�                                  �$EXTLOG_REQ        ��    �$EXTLOG_SIZ        ��    �$EXTSTKSIZ        ��  ��$EXTTOL      Dz  �A   �$EXT_BWD_SEL         �    �$EXT_DI_BWD S�������                  �$EXT_DI_STEP S�������                  �$E_STOP_DO        ��    �$FACTORY_TUN         d�    �$FDR_GRP 1T������  d 	                             	 YZ:���-�N#l�T.�E ��� ��� ��� 	                                      	 B���B�&uC�XB��EB�ArC��             	 A�)B[�B��DB�pA�w�B�             	 B/0�                                 	 ��@��%A%1A2����HAV�             	 A���B@��B$�A�]�A�׆B�             	 ��AW��.P����A �K���	             	 ?��A1��A�M{@��	A���A^�             
 F�4�B��DA�M{���HB:�                         c                 	 F?h FR� FR� Eu  Eu  D�               	 E�  E�p E�p D�  D�  DD               	 C�  C�  C�  B�  B�  B�               	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	 E�� E�� E�� E�� E�� E��              	 P]��P�W�P�W�M�DM�DK�y
             	 ?B�\?Y��?Y��?O\)?E�?0��             	 :I��:�o:�o9q,(9q,(9q,(             	 �s �n��M�{�ۦ��^.��]�             	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	  %U6 ��� ��� ��� ��� ��� ��� ��� ��� 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      
                                                                	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FEATURE U������   HandlingTool          �P��English Dictionary    ���Multi Language (GRMN) �)�`4D Standard           ��*Analog I/O            �	� Angle Shift           �Auto Software Update  �� �Automatic Backup      �â�Background Editing    �S
Camera I/F            ��c3CnrRndImp             �:AFCommon calib UIF      �2!�Condition Monitor     PiControl Reliable       �`Data Acquisition      B� �Diagnostic log        �h�Document Viewer       2��qDual Check Safety UIF ���sEnhanced User Frame   ����Ext. DIO Config       9�PKExtended Error Log    剟 Extended User Frames  �P&�External DI BWD       �L�FCTN Menu Save        �#�FTP Interface         ��Group Mask Exchange   �@`HTTP Proxy Svr        ���High-Speed Skip       ����Host Communications   G (Hour Meter            `�bI/O Interconnect 2    ���Incr Instruction      �?��KAREL Cmd. Language   4�BKAREL Run-Time Env    }�PKernel + Basic S/W    %�n�License Checker       A�LogBook(System)       ��TMACROs, Skip/Offset   4� MH Core               ���MechStop Protection   ��C�Mirror Shift          �ҀMixed logic           ����Mode Switch           4Zl4Motion Diag. Core     ��k`Motion Optm. Core     >`�@Motion Profiler       \��Motion logger         �h�@Multi-Tasking         �Sp�PCM function          I��|Position Registers    }0Print Function        ���Prog Num Selection    @ZpProgram Adjust        Nu��Program Shift         ��Z�Program Status        ��Program Viewer        �L�RDM Robot Discovery   �K�;Remote Conn Standard  �/�Robot Servo Code      ��SNPX basic            ���Shift Library          \�Shift and Mirror Lib   �D�Socket Messaging      �O �TCP Auto Set          �ZxTCP/IP Interface      4TMILIB Interface      �` &TP Firmware           �@.TP Menu Accounting    �$��TPTX                  -��Telnet Interface      ���Tool Offset           ��GTorque Simulator I/F  � �Touch Panel           ù!Trouble Diag. & Prev. �߯USB port on iPendant  Z��Unexcepted motn Check @�� User Frame            T�PVCalibration Common   ��RVision Core           �>�Vision Library        ����Vision SP CSUI        �K�bVision SP CSXC        ?�<Web Plus              s��Web Server            F�Web Svr Enhancements  ��iPendant              n�<iPendant Grid Display 2�iPendant Setup        ���4iRCalib. Standard     �  iRCalibration AAVM    ���Independent Axes      �� \Independent Axes      ¾�`Independent Axes      2�1�M-900iA/260L_iC       _8�Ascii Program Loader  ����Ascii Upload          �#�AutoMode TP operation &/� Basic Remote TCP      H��CE Mark               ����CPRUT                 8��CRT/Keyboard Manager  ��tCntrl stop by E-Stop  r�_�Collision Guard       ĩ~Collision Guard Pack  �^�Constant Path         �}�CornerDistance         p��Cycle Time Priority   �RDCS Joint Speed check +�`KDCS Safe I/O connect  c� �DHCP                  ��Domain Name Serv.     �9/Dyn Path Modifier     ��zEnhanced Dry Run      Q�O�Error Code Output     ���Ext Path Optimization  ��#Extended Axis Control d~External mode select  T�wPFRL Params            �f
�HMI Device (SNPX)     ���Integrated PMC        0�4�Internet Conn/Custo   �� Jnt Position output   9x�KAREL                 ��RMulti-Group Motion    �}8Operation logbook     �r�PC Interface          <��8PROFINET I/O          ��PROFINET Safety       ��ZPPROGRAM/JOG Override  >�P�Password Protection   � �PathSwitch            7 �SNTP Client           ���TCP SPEED OUTPUT      ���User Function          ��User Socket Msg       �~�VAG Package           ?:�VAG servogun setup    'L�VAG setup 3           ,�Y@Weaving               �<`�iRCalibration VAxis   ��Z64MB DRAM             �f�O64MB FROM             ���Arc Advisor           � �Aux Servo Code          �Cell I/O              �Common shell          r��Common shell core     |@30Common softpanel      ���Common style select    �xCorner Region         � UCycle time Opt.       U(�0DCS Pos./speed common �0@FDisp 2nd analog port  �0L�EMAIL Enhancements    � 0Email Client          �^�Enhanced Rob Serv Req  ��Enhanced T1 Mode      cxjpExt weave sch         ,�B,Extended Axis Speed   0�0Func stup             ;MC�OPT TP Ins            � PC Send Macros        }��Real Simple Syn.(RSS) q2@Requires CP           �PנRobot Library Setup   �&�Robot Service Request ���SMB Client            f`}SSPC error text       �P��Soft Limit            ���Space Check           ���TCP Speed Prediction  ����TCPP Extention        "V0Track Instruction     ? Tracking Softpart     bG`8VAG Software          ��histdpnl               F `�VAG V8.x Customizatio �>WVAG EMZ & EQ Tools    ^vRFREU late Updates     ���pUpdate VAG PMC        �SЩAscii Upload when arg rs�5Profinet and CD Setti ��"�*.pc protection and u �2��DryR.Skip PWF,VAGBCK  �&Activate CD Setting   � \�VAG Menu to Page 1    ��Implement Feedb.Tig/T ��'Fix upper limit of GO ���To fix skip problem   v���Files Updated          ��Activate CD-PS-Impr   �j�Diff.a.DryS.PN:FW-CHK ޚ�_Diff.a.DryS.PN:FW-CHK H�	CD:Fix SSTEP and BWD   ދFix.Er.after 8xVag_C. �@dUpdate several Issues U��Enh.Alloc.Mem.CD-Mot  ���To fix skip problem I �~Fix Err.Karel Var.Scr 08�<Fix DCS FB_CMP alarm  9�XFix overwr.VAG FUNC-M ܰ|�Restore Optimizations }�P0Fix.Karel User n.save ����ZIP cmd.er.handl.impr  ��yRestore Optimization  87� VAG Sign Off Function  #\�ATSHELL Heartbeat Opt ���No Outp.On/Off w.SRVO Ծ �Fix-PS strt move away ر��GunM.DO.Prot.Gen.Opt. �WFix iPend.scrn freeze ᰉ�P381+Investig.Patch   ����Fix ABC Over Run      ���Over.disp.unexp.clear  �PInv.probl.about PGPX  j�Res.TCPspdoutVar E-St 
8�Fix ABC Ov.load MSTP  r���Modification of iRCal  /�Unzip Inst+Improv.    �. Fix PGPX OX-144 probl LF�Enh.DryRunP.Canc/Res  8��Fix OS144 Motn-UserCa ����Improve VAG-Backup    �иImprove VAG-Backup    z���                      T4B��                      �@_�                      � 9�                      v��^�                      dâ��                      ``a �                      h�b��                      p���                      ��                      �r��                      H�k��                      �XvV�                      ��b�                       �^�                      l`�k�                      �U8�                      �p�,�                      *�p(�                      ��`��                      H����                      h�"�                      ޱ��                      ��a�                      ��*��                      ��Y��                      p�e��                      �}�n�                      �����                      �@�{�                      /P���                      ����                      ��H�                      �Py�                      G�!�                      �����                      �?@�                      �})�                      ����                      ���                      ����                      ���                      ǰ��                      n&��                      B L�                      "Y�P�                      ���                      ~˔�                      �iC�                      0���                      ;� �                      ����                      z��                      }` �                      ҙ^�                      R܎ �                      G �3�                      ����                       ����                      .^��                      ����                       �b��                      k� ��                      G U��                      ��9�                      � ]^�                      ���                      $�_X�                      w��                      |)��                      �}HP�                      �P��                      �`}�                      �\@�                      |�@�                      0}k`�                      aba��                      �J ��                      D@Kf�                      ߊ�.�                      qJa�                      OL�2�                      Nt�                      ��0�                      q ��                      �h��                      [p�t�                      @��                      �N���                      � H&�                      h P��                      Ww\��                      h`w�                      �C p�                      �� �                      (����                      ����                      ���                      b��                      4H��                      (8y �                       w|��                      �
�                      )�!�                      .����                      T=�@�                      ���                      P,,�                      N����                      2W��                      ˟ ��                      4.�,�                      �w<�                      ��W��                      }���                      ;^  �                      ����                      1}�[�                       :\�                      �4:�                      ���t�                      ��>�                      ����                      2����                       ,��                      ���                      H.���                      k\b��                      �cqb�                      rs�                      R��s�                      0w���                      ~�P��                      �Ə�                      {�}�                      Q��0�                      / <��                      UΒ�                      �
�                      +�}D�                      P��!�                      ����                      ����                      v��                      k��                      �"}��                      �~���                      �v���                      ����                      �؁}�                      2r���                      �2��                      �:��                      �f��                      �<�A�                      W���                      ��x~�                      ��X�                      Z9W�                      PK~��                      �n�;�                      ��T�                      ePZd�                      Y�B��                      �~��                      �����                      ��9�                      �����                      ��t�                       ��q�                      $����                      B���                      Ò��                      ���8�                      �����                      r��                      ����                      �
���                      � .�                      $����                      �+�                      �d��                      :�[��                      P9�                      *�y��                      a
��                      EA��                      0Bj��                      bs��                      ~���                      ����                      O�A��                      �� �                      ��0`�                      ~���                      ����                      F�`�                      !��                      $@PP�                      ��B��                      h`�                      �H-�                      n@��                      �9%��                      "4���                      툞g�                      ��`��                      �uD��                      ���8�                      ��M��                      ���                      ڥ6P�                      ��8�                      y�.�                      �I 
�                      >Q΀�                         �                      ?�� �                      ���(�                      ƥ�>�                      ����                      P��                      ����                      � X�                      �Qf!�                      Y�r�                      �$�                      $�B��                      �(�                      �?b�                      `�d�                      }k)U�                      �� d�                      }
`��                      ���!�                      JX���                      ?�u��                      ��B�                      @�l�                      �0�?�                      `X��                      @D�                      �����                      ��1�                      �����                      ��T8�                      ��#�                      �����                      �H�                      �*�                      ��_|�                      �-*�                      ^p�                      ���                      ��t�                      H��0�                      �r�z�                      ���8�                      (� h�                      �@8��                      w��@�                       A� �                      ��8��                      ��o��                      �|c:�                      �Bԃ�                      �d �                      ����                      2�`�                      ?�C�                      ��Y(�                      �h��                      ��                      �r�                      �0���                      ����                      ʢ�`�                      a� ��                      �����                      ���a�                      ��Cp�                      rq �                      r���                      �@��                      ���p�                      ��	��                      ��                      ��D�                      r� �  H552  h$�H521   �}H532   �R782     H550  8~FJ614  �EԾATUP  U>J545  �w�JJ616  ��Y�VCAM  ���CRIM  �U�CUIF  t�� J628  ���6CNRE  �@R631  �@RSCH  ���DOCV  "O DCSU  �<@�J604  1���EIOC  `8�R542  �� �R696  �r�7ESET  
���J516  ���mJ716  ���MASK  ��$�PRXY  ��I�J627  �@��HOCO  q(�J513  ���J542  �� J510  ���$J650  �K�J539  ��HH510   ;��LCHK  �@OPLG  z��J503  s�HMHCR  �� MCSP  �x�FJ506  ���J554  � ?�MDSW  ]��MDCO  �x� OPCO  R��MPRO  ,�m�R637  ��J600  ���PCMF  �,�J514  t��fJ507  ����J515  |��J517  �+�@J505  ���PRST  Ł� J697  � ��FRDM  ���RMCN  ؁�H930  �Z@BSNBA  T��=SHLB  ���SMLB  � R636  �~� J520  ���HTCP  � $TMIL  0(�0R789  &0X*TPAC  �� �TPTX  B�0TELN  0�J509  �0�J882  0�/0R781  K0�?J958  L[0�J957  �0�\UECK  �1�UFRM  j�� VCCM  �OH VCOR  (��VIPL  K[��CSUI  ��PCSXC  �KG�WEBP  0:E�HTTP  � 
�R626  �FO CGTP  \MOIGUI  �@�IPGS  A�' IRCL  ±��J888  P?@4H895  P"�H895  _�_~H895  �K�FH621  ���-R796  �{|R507  N�  J698  �0 R657  x���J618  Q��J858  �� DJ535  �� J570  �d0�R534  �o`RJ684  � ~R663  �x��R748  ��JpJ523  ��pJ555  q�|�J568  ���R526  _��J755  ��8R739  <ѧJ985  t~��J527   ���J829  ��d8J518  �9�J569   �LR651   �BR553  \��?J760  J`$R558  TmJ966  x�,�R632  ��S#J601  �0�J695  ���R641  �vNJ930  ���~J931  ��^ J579  ��L�J541  ����J693  ��8�R610  iT�J694  ���|J986  ��} R648  ��J658  0�"�J653  � <�J656  �@�J504  5 J996  �4D064  ,^�F064  ɡ �R666  ���SVMO  `�MCLIO  }��R645  � hCMSC  |�ЂCMSP  � PfSTYL  �|�R654  8�CTOP  ��TDCSC  h��R528  ��}JNN8  ��JNN7  `� 6ORSR  �hL�R680  ���J881  � $�EXTS  |�s�FCSP   �VOPIS  |��SEND  ߠ�R679  B���CPRQ  J nRLCM  Hm��SRSR  �b�R677  ϩ}ETSS  G��~SLMT  }�Y�J609  �JaJ524  p�nTCPE  �+��TOAW  ��TRAK  �K#FVAG    �IPNL  ���VAG1  �08EZEQ  �}��UPD3  ?��HPMC3  ��� P137  b�iE001  �P�E002  �x�E003  ��a E004  XM��E005  ���E006  ��P170  H � P171  DfvE007  t�� RT22  C2�E008  ���E009  @1�P208  8�@�E010  � 8rE011  ��a RT23  �@��P213  ��PP225  ��"P230  ~:�P231  8�� E013  �bP238  ��2P244  �a�E014  �� �P246  k��S300  �`�P275  f�?P276  �a 0E015  ��H�P381  k�*�P477  f�~P501  8ࡄP525  ����P537  r���P333  p.�E016  �2��P307  b<�P576  l��P604  �T~E018   D��P623  { ÂF001  1� �F002  z$��      �����      <����      �~��      <��      �0qH�      ���      0���      �<�9�      �4��      �2���      Hak��      �� �      ,����      V!���      ��a�      4&��      ~֐P�      ��@��      ޠX~�      �X�b�      �B��      ����      ak �      �^ ��      �`���      �1ց�      |0��      }�J@�      0��0�      �'�      �6���      �~h�      @��`�      ����      K7���      ����      �/�      �^�Q�      ��h��      ����      X�� �      � r�      ����      ��=��      v�{ �      ��¥�      j0?�       ,*o�      �+ �      �b  �      o���      J @Z�      o��X�      ��o"�      bZ1��       �ނ�      iC L�      �o�      oP�#�      l$0��      ���n�      ~����      HX�      ����      � Ц�      瀙a�      �A~��      � J�      ����      �ut�      H��^�      ���J�      [�Ћ�      4,��      ��q8�      �k�b�      �����       ���      �  ��      �QP�      ����      ~_��      @!��      ��:1�      ,|��      � ħ�      �@_ �      ���      ����       CK��      �B� �      }JJ��      Pp���      T���      ؅��      :���      �s��      N���      � >�      �H��      (�Ѧ�      ��{8�      � �      �A���      Hbs�       Ժ��      ��H�      �V��      E���      �x���      !��      :���      ���0�      � ���      ��H�      R����      `�X�      �Ђq�      0���      9]0 �      %��      �J��      К���      w��      ��e�      ���      r�j �      {��q�      ����      H�L�      �T��      =\��      `��      �j� �      f�;��       ��      ��{�      �?���      ���q�      G����      �����      ����      �\��      @(.��      ���H�      &� ��      ����      ��~�      ?�8�      8�`�      0~jF�      TP��      � �n�      ���      >,"�      PQ�      �T��      ��̲�      x2,|�        B0�      �j2C�      �[0�       ,���      J� ��      ��[�      mk8��      `(���      �� ��      �b0�      �� ��       4T��      ���/�      �zT�      �4���      ����      �B��      �?~�      �!��      0! 0�      _*_p�      XL�E�      P�wP�      �P���      �_�V�      PD�R�      ��F��      0��_�      Ҝ�L�      ���      ����      X���      pNT��      ��~��      �r��      �?��      �����      ����      T��h�      �`~}�      a���      �\�      �NTH�      8��H�      t~�&�       �K�      ��o`�      �����      �Db��      �2��      ���0�      �D�       h��      ��\�      t��      � ��      n�r�      ����       ���      < ��      �~ �      �`@��      ����      �8z�      IRT�      �iq��      ����      X��L�      M?���      $S��      @
�9�      >�C�      �����      Zޖ��      A���      �����      ����      ���      �m�^�      �A�      �� �      B၌�       ���      Ѭ (�      �v��      ߠ���      ��      ��V��      ����      �"�4�      O�Z��      w�V��      �r���      ��L�      �9 `�      ����      9l�w�      Hm� �      ����      �J`T�      Q�$ �      l���        ���      �� &�      �� ��      ��~r�      ,�`��      �:��      f�!��      W
Ě�       ���       ���      �r��      �_�      J!>R�      �� �      Q����      ~rߏ�      �T�A�      ~�4�      2�P��      Д:��      �F}x�      ��4�      �  �      ��      4`�      ����      �_?  H552      :�� H552       HH552      �Ѐ�H552      �8��H552      <��H552      w�H552      ҀXH552      X$�/H552      �R2/H552      �l�H552       ��H552      } �0H552      ;�  H552      ��0�H552      ?B�H552      ��#H552      9 0H552      ||yH552      �pH552       
8�H552      9 ? H552      ���H552      `�� H552      D ��H552      }HH552      ] \�H552      @|SH552      ��@H552      9J H552      ���H552      P	D_H552      Q;~H552      @��lH552      �F!H552      dx�>H552      j�PH552      �X(H552      |�H552      r}�H552      �8� H552      �}EH552      P_�UH552      
l|�H552      Ш�"H552      �ev`H552      &Q?`H552      0[$PH552      ��JkH552      aC@H552      ���}H552      �i}�H552      `})�H552      v��H552       �bH552      �QH552      
&pH552      j`}kH552      ���H552      q�H552      �ԐH552      ��H552      -���H552      `PVH552      ,���H552      PK�FH552      {�A�H552      <ƍ�H552      A��H552      X�(H552      �h H552      }�@,H552      \|	�H552      (?�H552      
(�H552      ���iH552      $��H552      ���0H552      7�� H552      E(Z�H552      qj�}H552      낿�H552       ��H552      ��l�H552      ��6H552      G+1�H552      f0�H552      ���|H552      ����H552      �^�H552       �H552      ��	JH552      ,�}�H552      �0�aH552      =@ H552       L8aH552      @�1�H552      �$�H552      �.]H552      � u5H552      �V�H552      �@�H552      7���H552      ���H552      �ӰH552      },.@H552      AH552      ��.H552      i{l�H552      ; �H552      � �8H552      l�H552        �H552      T�6�H552      ���H552      ��|�H552      0~�H552      �kH552       ���H552      ~ �H552      \�RH552      ���TH552      D���H552      odH552      f�ZH552      �b�H552      �8?H552      �@�aH552      0"vH552      �H552      yD��H552      ��~�H552      ���H552       b��H552      � @�H552       �<H552      ^��PH552      b�H552      Ќ��H552      ���H552      �baH552       a� H552      �bbH552      =rbH552      �2H552      Q sH552      8z0H552      �8� H552      ^2�H552      ���H552      �t� H552      �t��H552      ����H552      �@�H552      8�H552      ���H552      6���H552      ���H552      �`�hH552      �*~6H552      ����H552      ����H552      ��ؐH552      {h$�H552      }��H552      _;kH552       �H552      `[ H552      � x H552      �g�>H552      ��@�H552      �H552      �JH552      �� H552      䒠�H552      �d�H552      p"�b           ��<           �BaN           �B           \~�           �b�           ~��)           �ZB           ��           1��|           P�           X��           ��X           ?8}�           ����           ����           �Z           ���M           �RL�           o��            � �1           D�
H           � @           �Hvd           ��)�           ���           ��(           ���           h$��           �1;           �9?�            ��           ���           |�b           �Q6            �+�`           B�T�           ��`�           ��           j�8           �V�           �c�           ���|           x���           $�R�           h��            ��           $�            A���          �M@�          �*��          А���          l ���          �Ɯ��          �`$��          ����          <����          �h���          � ] �          Y6a^�          /A���          ����          ~��          a*��          *~�>�          ~�d��          ���w�          �aA�          �p�;�          T���          �i�          |��          8��v�          ���          1�0��          K���          ��|�          8P�`�          ��a�          ���          �F��          � ��          �
���          �`�          `Q� �          $@;P�          � �P�           |Z��            ��             �          �<�          <���          �@��          �a �          �� ��          ɡ (�          ���h�          |;�M�           �h�          ����          ~P���          |X �          ��B�           |�          }�>��          �<�          �Eh�          6� }�          Z�K��           &��          �@��          �B��           ��          ��k�          ��h��          { ��          �Yֱ�          ��0��          �ؾ�          C���          �X�          ?���          ��}J�          �P�k�          ѐ�          }����           ���          � �          ? X|�          |oeI�          �,�          �Ё�          �l��          s�0�          ����          ��J2�          B����          Ir"�          ~���          A W�          L��          �d|
�          Ҍ0��          Щ^��          J ��          �1�|�          }��@�          ��,��          (f�,�          �����          �s�H�          ����          y�[�          �t��          � ���          ?�<�          �����           0���          P���          
@��          ���}�          (��          ��p��          �K$�          �4���          "��          J��I�          �K8��          �@H�          2 +�          �B���          � D*�          ���H�          >�F�          B���          _��          ��          N`�          �w��          G=���          r���          ����          �*�K�          /<�V�          ��~��          ����          �� ��          �����          ���`�          � hy�          �5���          ��-�          ��(��          �����          �� �          �;�(�          �8���          $��          /0�y�          ��@��          E�@��          瀃�          :�?�          P�� �          U��          ����          �����          �W���          �����          � b�          ��(��           DN��          "����          �jVP�          ����          �U���          �Q
�          UV�0�          ����          KK���          X@ߑ�          �@'�          O\_��          �pF�            R�          ���          �~���          ����          ��\}�          ��          _��[�          �*��          �T��          ��A��          �20�          z��'�          P�          ��a9�          DW��          ���r�          p�C�          �pL��          �G�p�          �Xj��          �����          �ޏ��          0"�Q�          t�p4�          x�p|�          z��          ®��          Sɲ��          ��"�          n���          �!�R�          RM.��          όϞ�          ��(��          a � �          �+���          Z����          ����          ]'��          �����          x,
�          �z�0�          �h��          �|x�          ��� �          O�:�          �d��          �g��          b�-�          pT���          X��\�          ��o��          ��v�          �����           e��          (̃�          �;/��          ����          6Ȳ��          JY@�          CI�          �R_d�          HLM�          �&�          �jH �          "5�x�           PL�          "_4X�          �/�B�          ?8�          H�          o���          HJ�          J# ��          Q�9{�          0}k`�          |�Q�          3`Y�          |e4�          A� �          e�          �N}�          ��LP�          �T��          �?�l�          ����          A� �          �00
�          �0m<�          �݁�          l�g��          ����          �c���          �zѠ�          ;�� �          �YH�          � ��          �Pp��          �|l[�          ��S�          U$� �          OHG�          bQ���          ����          ���          Z���          x���          �� �          $��          � ��           ����          ��_�          B �D  STD   ��X�LANG  ���LANG  ��� STD   ���STD   ��ASTD   Y.�eSTD   TzюSTD   4��STD   }kSTD   9> �STD   �~��STD   �)LQSTD   ����STD    � STD      STD    ��STD   ;��STD   ��\�STD    7�STD    �b/STD   "�HSTD   (�STD   ���STD   (�l STD   � 0STD   �);�STD   #� 8STD   �@`STD    �  STD   X @STD   <<JSTD   2@(STD   k1LSTD   � �STD   ! 0NSTD   	��STD   �H�STD   �/STD   �0�STD   4m�STD   � �STD   �0��STD   ���STD   �f�STD     STD   A��OSTD   KX �STD   �@k�STD    ���STD   ��HSTD   8��STD   ��}STD   |�0STD   � hSTD   }�4STD   �O�CSTD   ��B�STD   �STD   �_STD   ��x�STD   �_�STD   K�� STD   �P0�STD   ��STD   C�_STD   CB`�STD   f�T@STD   !�{STD   �I�JSTD   o�TESTD   �C�`STD   dE�STD   E�"STD   	<R STD   ��STD   ����STD   ��� STD   w�}STD   �dESTD    &RSTD   �� "STD   �� STD   ;��PSTD   <�?!STD   �A�STD   @�H STD   ��X STD   ���STD   $�|�STD   ���GRBT   A��RBT   i��RBT   �⁑RBT   �~ �OPTN  br�0OPTN  �PqiOPTN  "d!OPTN  s<��OPTN  @�DOPTN  D�frOPTN  �$�COPTN  �XG�OPTN  �A)OPTN  ���oOPTN  ���OPTN  M� �OPTN  "� $OPTN  �a*�OPTN  ~��OPTN  _�(OPTN  ����OPTN  =R��OPTN  a|sZOPTN  ,�OPTN  f��POPTN  �rFOPTN  R,v4OPTN  ^��jOPTN  �p�AOPTN  &\q�OPTN  6�H�OPTN  @�pcOPTN  O���OPTN  �7@OPTN  @= OPTN  �AG�OPTN  +��OPTN  �O��OPTN  �+!_OPTN  �Ƀ�OPTN  �h�OPTN  0�d@OPTN  7�~�OPTN  �`OPTN  ���$OPTN  �L`OPTN  �<��OPTN  x�!�OPTN  ���OPTN  J(�DPND   }@rDPND  1A�DPND  �@��DPND  0��HDPND  �L"ODPND  ��NADPND  az mDPND  �8�@DPND  k�@;DPND  ��RDPND  ���DPND  ��p�DPND  &ڝ�DPND  �xHDPND  8���DPND  � rDPND  N�UDPND  �A?DPND  W]�DPND  G��DPND  �
��DPND  ����DPND  �DPND  �� rDPND  ^�;�DPND  D"DPND  �/DPND  �,DPND  ���DPND  �N�DPND  ����DPND  �� (DPND  ���/DPND  u0��DPND  ���DPND  ( 8CUST  �FCUST   @�PCUST  O?��CUST  HrfCUST  �8Q`CUST   hLCUST  ���CUST  pK?�CUST   TzCUST    �CUST  ���CUST  .parCUST  �)p�CUST  mal-CUST   >- CUST  N)orCUST  PaPCUST  �N CUST  INPUCUST  z�)RCUST  �/�&CUST  C�@�CUST  d hfCUST  Pln@CUST  End)CUST  022ACUST  UninCUST  0 r%CUST  co�CUST  �`CUST  �4� CUST  8p)CUST  an�@CUST  '�3CUST  BFCUST  V>)pCUST  5�F	CUST  *2qCUST   tf_CUST  o2CUST  g�pCUST  ilZpCUST  Xp�CCUST  0�qXCUST  C�1 CUST  !�O�CUST  p�rnCUST  eGc)�      N^e�      2��      :np �      1F	v�      radi�      �_�_�      V���      +)&�      |m�      �=oO�      o_Kc�      A�~�      � ��      I�Iu�      L�I�      umb�      �N1,�      "�G�       �C��      �zDr�      � E��      eck_�      D02�      �IsN�      able�      �{2_�      pcon�      ntk��      ыn��      �@SH�      Pd�_�      ~0(�      ;��3�      6.4��      dsb��      �0hc�      
 ��      AR�T�      �OMO�      E ���      P:0a�      ��0�      �p{��      @ex�      >��D�       �2��       �B>�      del��      @R2�      D��[�      H+�      @2�M�      �4� �      ���       f p�      ͱF�      o��      Am���      �р#�      �2�      0#��      ���      inp�      ����      6�nd�      �NIS�      potT�      andl�      Disp�      rc���      �Ro/�      �l���      E�Q��      ��E�      �# �      %x((�      �POS�      ��$%�       �      gr��      SpNo�      e_
��      nPͰ�      t1:�      �AO��      @p�q�      wp���      =�TE�       :���      axis�      mt��      I� �      ��'��      lrnm�       [cp�      prv�      ���O�      Yo���      ��]��      p��      �r���      Clo��      |��      ouك�      �ЀM�      B� �      4�A �      � � �       @@��      �o9�      �~@�      �k ��      k9A�       ���      �P0}�       ?A��      ���      � ���      �� ��      >��J�      J� ��      �� )�      �P<�      �8C�      J�9�      ov�      `��      ƒ8�      �� �      ���      �� �      �� 
�      ?�� �       ��      w��      sol��      �dec�      %pe�       t1_�      f �u�      �b{c�      �oCi�      0�t��      ҭq8�      s'�1�      Pp���      Delt�      �n���      l��w�      ����      in�      to_g�      vrĵ�      � _�      t¡��      q����      ��_��      Կ���      =Rr��      �9���      aա��      e-p��      r�`��      ώ�0�      jb���      :  ��      �CPl�      X�m)�      �����      o6��      ����      � �n�      �fil�       �U��      �1�`�      _&���      ���      ����      ����      mp_m�      �va��      �irr�      �Z�      ��R�      S�j��      :� E�      es2w�      n�l��      �`er�      c�l�      5f),�      � R��      �g� �      ��	�      v�-d�      	 f��      X�D�      Tool�      � fr�      �� o�      alw!�      �����      h� %�      �G1�      J߰\�      S q-�      rgi)�      ���p�      �X��      MODE�      E�`��      =�H��      u8��      oa��      '3: �      $�$�      =4  �      �A)�      � ���      5�/4�      Pp.�      �E���      �0��      dY���      -R�P�      �f �      �`���      � OP�      r1�?�      0)O�      �O�O�      �O�O�      l�?x�      ldC_�      B,pO�      O�_��      Mark�      cXoj�      xGq=�      b L�      � $��       O�'�      .t6j�      h��      ���f�       a���      �GrC�      + A��      y�Wo�      `aAr�      �p_��       �� �       REP�      $FLA�      �Fp5�      ?NIS�      low��      ����      ����      Ï��      �����      ��SW�      �KED�      NORS�      �T���      L�$�      B�T��      ��OG�      �Ȧ��      �>��      C�E�      <����      �Կv�      Ͽ1�       FIL�      ��W��      �Ϛ��      �����      �H� �      ����      �ȯ�      � f��      (����      ���&�      1���      K����      3)99     ����$FEAT_DEMO U������   �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                            �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �            �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �                �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �$FEAT_DEMOIN         ��   �$FEAT_INDEX         ��   ��$FILECOMP V�������        �$FILESETUP2 W�������  �  N   N �$FILE_AP2BCK 1X������  �)MAKRO900.TP                               %MAKRO900                                 %MAKRO900                                  )MAKRO910.TP                               %MAKRO910                                 %MAKRO910                                  )MAKRO920.TP                               %MAKRO920                                 %MAKRO920                                  )MAKRO930.TP                               %MAKRO930                                 %MAKRO930                                  )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_APPBCK 1X������ 2 �)*.VR                                      %*                                         %                                           )*.PC                                      %FR6:*.PC                                 %                                           )*.TX                                      %FR6:*.TX                                 %                                           )*.FVR                                     %	FR6:*.FVR                                %                                           )*.STM .STM                                %FR:*.STM .STM                            %iPendant Panel                            )*.HTM                                     %FR:*.HTM                                 %                                           )*.GIF                                     %FR:*.GIF                                 %                                           )*.JPG                                     %FR:*.JPG                                 %                                           )*.JS                                      %FR:*.JS                                  %
JavaScript                                )*.CSS                                     %FR:*.CSS                                 %Cascading Style Sheets                    )
ARGNAME.DT                                %FR:\ARGNAME.DT                           %ARGNAME                                   )	PANEL1.DT                                 %FR:PANEL1.DT                             %iPendant Panel                            )	PANEL2.DT                                 %FR:PANEL2.DT                             %iPendant Panel                            )	PANEL3.DT                                 %FR:PANEL3.DT                             %iPendant Panel                            )	PANEL4.DT                                 %FR:PANEL4.DT                             %iPendant Panel                            )SHELL.VR                                  %SHELL                                     %�                                          )ZG_MENUE.VR                               %ZG_MENUE                                  %�                                          )
EINGABE.VR                                %EINGABE                                   %�                                          )SUMM_VAG.DG                               %FR:SUMM_VAG.DG                           %�                                          )TPE_STAT.VR                               %TPE_STAT                                  %�                                          )	IO_SET.DT                                 %FR:\IO_SET.DT                            %�                                          )VWEMZROU.VR                               %VWEMZROU                                  %�                                          )VAGBCKUP.VR                               %VAGBCKUP                                  %�                                          )
TPEINS.XML                                %FR:\TPEINS.XML                           %Custom Toolbar                            )PASSWORD.DT                               %FRS:\PASSWORD.DT                         %Password Config                           )VAGCONF1.XML                              %FR:\VAGCONF1.XML                         %�                                          )EXTSERVO.VR                               %EXTSERVO                                  %�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_DGBCK 1X������ ( �)
SUMMARY.DG                                %MD:SUMMARY.DG                            %Diag Summary                              )
CONSLOG.DG                                %MD:CONSLOG.DG                            %Console log                               )	TPACCN.DG                                 %	TPACCN.DG                                %TP Accounting                             )FR6:IPKDMP.ZIP                            %
IPKDMP.ZIP                               %TP Exception                              )MD:MEMCHECK.DG                            %MD:SUMMARY.DG                            %Memory Data                            �)MD:SHADOW.DG                              %MD:SUMMARY.DG                            %Shadow Changes                        �g)	FTPLOG.DG                                 %MD:SUMMARY.DG                           %Comment TBD                           \+�)ETHERNET.DG                               %MD:ETHERNET.DG                           %Ethernet Configuration                    )MD:DCSVRFY.DG                             %MD:SUMMARY.DG                           %DCS verify all                        �z�)MD:DCSDIFF.DG                             %MD:SUMMARY.DG                           %DCS verify diff                       �z�)MD:DCSCHGD1.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �O,)MD:DCSCHGD2.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �O,)MD:DCSCHGD3.DG                            %MD:SUMMARY.DG                           %DCS verify diff                       �O,)UPDATES.DAT                               %FRS:\UPDATES.DAT                         %Updates List                              )
PSRBWLD.CM                                %FRS:\PSRBWLD.CM                          %PS_ROBOWELD                               )MD:SMTPLOG.DG                             %MD:SUMMARY.DG                            %SMTP/Email diag                       �-�)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_FRSPRT  �������    �$FILE_MDONLY 1X������    
 �)�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FILE_VISBCK 1X������ 
 �)*.VD                                      %FR:\VISION\DATA\*.VD                     %Vision VD file                            )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          )�                                          %�                                      ��%�                                          �$FMR2_GRP 1Y������� �C4  B�   	                             	 E�� E�� E�� E�� E�� E��              	 P]��P�W�P�W�M�DM�DK�y
             	 ?B�\?Y��?Y��?O\)?E�?0��             	 :I��:�o:�o9q,(9q,(9q,(             	 A�  A�  A�  A�  A�  A�  A�  A�  A�  BH   	 C�  C�  C�  B�  B�  B�                  	 D      CH          Da               	 @UUU@UUU@UUU@UUU@UUU@UUU             	                                      	                                      	 :�}:��:Bj9���9�f,9֯�             	                                      	                                      	 F?h FR� FR� Eu  Eu  D�               	 E�  E�p E�p D�  D�  DD              C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     C4  B�   	                             	                                      	                                      	                                      	                                      	 A�  A�  A�  A�  A�  A�  A�  A�  A�       	                                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$FMR_CFG Z������� T                                                                                    �$FNO �������F174554               �$FRM_CHKTYP  ����   ������$FROMCHK_MIN        ���  X�$FSSB_CFG [������                                                                           �$FTP_DEF_OW         �    �$FTP_DIRCOMP         �    �$FUNC_SETUP  �������                                                                                  �$GENOVRD_DO        �   �    �$GENOVRD_THR         d   �   d�$GENOV_ENB         �   �$GRAVC_GRP 1\������  �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            �    	                                          	                                          	                    	                            ��$GROUP 1b�������                       8�?�              ?�              ?�                  8��;�.�   ?�  �   ?�  �   ��  �   �;�.ĕ�3�&ffCe33    C�  CH                                                             Cx:�               B�                                                                 8!�?�              ?�              ?�                  8!�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   81�?�              ?�              ?�                  81�?�              ?�              ?�                  C�  C�                                                              �                  B�                                                                   8A�?�              ?�              ?�                  8A�?�              ?�              ?�                  C�  C�                                                              �                  B�                                             �$GRSMT_GRP 1c�������      C�      C�      C�      C�  �$HOSTC_CFG 1d������ ��                  	FTP       �            �                          172.26.26.230                e                                                                                                       e�                                                                                                      172.26.26.230         e	cfg_fanuc                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e	anonymous                                                                                                         �$HOSTENT 1e�������  P!�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !�                                        !�                                  !QUICC0                                  !172.26.26.84                      !QUICC1                                  !�                                  !QUICC2                                  !�                                  !ROUTER                                  !172.26.26.1                       !PCJOG                                   !192.168.0.100                     !CAMPRT                                  !192.168.1.10                      !CAMRTR                                  !192.168.1.10                      �$HOSTNAME !�������!KJLTVL111120R01RS--KU1            �$HOSTS_CFG 1d������ �Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  Auto-started      	FTP       �            �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                                     	SM                     �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                            �    �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �                  	�          �             �                          �                             e�                                                                                                      e�                                                                                                      �                      e�                                                                                                                  �$HOST_ERR f�������                    �$HOST_PDUSIZ     ^  ��  >�$HOST_PWRD ?������   �  backup        guest         guest         guest         guest         guest         guest         guest         �$HSCDMNGRP 2g������� �      d               K       	P01.04 8   	   E  
  �  ?  �  �             	 ���������������������X             	   ;  �  U  
  
+  	             	 �������3����������������             	   �  b  �  h  �  {             	 ���	�������������\���             	   �  �  �  �  q                 d 	   E  
  �  ?  �  �             	 ���������������������X                  d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                           d               K       	12345678   	                                      	                                      	                                      	                                      	                                      	                                      	                                        d 	                                      	                                     �$HSCD_GROUP 2h������      	HSCD01.02         �                  �                  �              �$HSCD_QUPD         �   �$HSCD_UPDTYP  �������   �$HTTP_AUTH 1i�������  <!iPendant                          �                    !KAREL:*                           �                    !KCL:*                             �                    !VISION SETUP                      �                    !�                                  �                    !�                                  �                    !�                                  �                    !�                                  �                    �$HTTP_CTRL j�������                 
 ��FFF9E3                       FRS:DEFAULT               FANUC Web Server             
�$HTTP_PWRD ?������   �  �              �              �              �              �              �              �              �              �$HWR_CONFIG k�������  f                    �$IBGN_CFG l�������       2   @   <#�
<#�
<#�
BH  <#�
<#�
<#�
CH            4   <#�
        �$IBGN_DEV       ���   �$IBGN_ERRIO m�������                �$IBGN_EXDAT n������   �            �$IBGN_EXFLG            �    �$IBGN_FIL o�������                    �$IBGN_FTP p�������                    �  �	MERCATOR  	RECORD    	R_ACHS    	R_ISTW    IBGN  IBG   	SENSPS    TXT   999   	Keine 0                                     %IBSCRECS                               8�%IBSCRECE                               ��           �$IBGN_LMTN  �������                 !                                                                                                        �$IBGN_SBADR      ���   ��^�x�$IDL_CPU_PCT      B�   B��$IDL_MIN_PCT      B�   =gF��$IGNR_IOERR        ���   �$INPT_SIM_DO        ��    �$INTPMODNTOL         ��    �$INTP_PRTY        ��    �$IOLNK 1q�������                                                                                                                                  �$IOMASTER         �    �$IOSLAVE r�������    �$IO_AUTO_CFG         �    �$IO_AUTO_UOP         �    �$IO_CYCLE         �    �$IO_DEF_ASG 1s�������              d                     d                �   c                �   c                  
   c                  
   c                                                                                                                                                                                                                                                                                                                                                                                                                 �$IO_DEF_NUM     ����   �$IO_IPCHE         �   �$IO_RTRY_CNT      ����    �$IO_SCRN_UPD        ��    �$IO_UOP_CFG t�������    �������������������������$ISDT_ISOLC  �������                  �$J23_DSP_ENB  �����������$JOBPROC_ENB         �    �$JOG_GROUP 1u������� 8   d8�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8!�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d81�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                   d8A�?�              ?�              ?�                  ?           �                  �                  Q�                                                                                  Q�                                                                                                                �$JOG_IN_AUTO      ����    �$JPOSREC_ENB         �    �$KANJI_MASK        ���    �$KAREL_CFG v�������          �$KAREL_ENB         �   �$KCL_LIN_NUM         �   �$KEYLOGGING  ����   d�   �$LANGUAGE �������ENGLISH       �$LGCFG w�������         ��   x  �  �  H  �   '0           �                     MC:\RSCH\00\                 �$LN_DISP x�������                                                    �$LOCTOL      Dz  �A   �$LOGBOOK y�������   d               d  X                                                                                                                                              	LOGBOOK            ��                                                �$LOG_BUFF 1z�������                    d                         d                                                                                                                                                                                                                                                                                                                                                                                   �$LOG_DCS |�������    =���                                        �������������������������������������������������������������$LOG_DIO 1}�������  ������������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ���������������������  ����������������������$LOG_ER_ITM  ������� d                                                                                                                                                                                                                                                                                                                                                                                                                 �$LOG_ER_SEV  �������   �$LOG_ER_TYP  �������                                                                                  �$LOG_REC_RST         �   �$LOG_SCRN_FL 1~�������    �                                                                                                                                                           �$LOG_TPKEY  �������                 �$LONGNAM_ENB         �   �$LUPS_DIGIT         �   �$LU_LOADPROG %�������%UP024                                 �$MAXUALRMNUM       ��   
�$MAX_DIG_PRT        �   �$MCSP ������                               d                �$MCSP_GRP 2�������  �   2     	   �  q  �                         	                                      	                                             	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                              	                                      	                                      	                                              	                                      	                                     �$MD_LDXDISAB  �����������$MEMO_APNAME ?������� 
 �              �              �              �              �              �              �              �              �              �              �$MISC 1��������  � 	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                          	                                      	                    	                    	                                      	                                         �$MISC_MSTR ��������    �$MISC_SCD 1�������� 
 � 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                     �$MKCFG ��������                       �$MLTARM_CFG �������          �����������������������������$MLT_GRP_DO ��������         ��L��                                                                                                                                        �$MMETPU       ���    �$MNDSP_CMNT         �   �$MNDSP_MST ��������                                              �$MNDSP_POSCF         �   �$MNDSP_PRPMT         �   �$MNDSP_PSTOL 1��������  4@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
@   <#�
<#�
 	 <#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�$MNSING_CHK         �    �$MODAQ_CFG ��������                             �$MODAQ_DEV 	�������	MC:       �$MODAQ_HSIZE  �������   ��$MODAQ_TASK %�������%$123456789 123456789 123456789 123456  �$MODAQ_TRIG 1��������  l������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ���������������%�                                      ������%�                                      ����������$MODAQ_TYPE      ����   �$MODEM_INF 1������� `)AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          )AT&FV0E0                                  )AT&FE0V1&A3&B1&D2&S0&C1S0=0               )ATZ                                       )ATH                                       )�                                          )ATA                                       )�                                          )�                                          �$MONITOR_MSG ?	�������   	EXEC1     	EXEC2     	EXEC3     	EXEC4     	EXEC5     	EXEC6     	EXEC7     	EXEC8     	EXEC9     	EXEC10    	EXEC11    	EXEC12    	EXEC13    	EXEC14    	EXEC15    	EXEC16    	EXEC17    	EXEC18    	EXEC19    	EXEC20    	EXEC21    	EXEC22    	EXEC23    	EXEC24    	EXEC25    	EXEC26    	EXEC27    	EXEC28    	EXEC29    	EXEC30    	EXEC31    	EXEC32    �$MOR_GRP_SV 1�������  ( 	 ?�
��
�?
�4�2���9���             	 B�                                  	 B�                                  	                                     �$MOTASK_DATA  �������    �$MPL_NAME !�������!Default Personality (from FD)     �$MRR2_GRP 1����  	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                                
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                   E�  E� Fp          	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$MRR_GRP 1�������  `    X, �    �� @D�  D�  ?�  ?�  X,?   ?�      @_f�D�  D�                             ;�	l?�   	 ���T��    	 �^� � � � � � � 	 K�s�K�ԼK�@K�@Kv(�KK             	                      	   �  �  �  �  �  �  �  �  � 	 ?�f�?�?�;g@
�@
�@_f�                     	 �Iۿ��6�ws�����X���             	 �4    ��Pô  ��  ô               	     >LU!���]    ��6X                 	                      �   �   � 	                                  	   �  �  �  �  F  m  �  �  � 	                                      	  	'� �  �  I� �  ��             	 :�È:�È:�È:�È:�È:�È=���=���=��� 	  @ @ @ @ @ @             	   �  �  �  �  �  �              �    	                                	   ��  ��  ��  ��  ��  ��  ��  ��  �� 	 @I�?��6?��@��@�X@��             	 C4  B�  B�  C�  B�  C�                 �C�   	 �#����       	        � � I       	 C   C   C   B   B   B                 @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  I� �  ��            �   � :=              �  @?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	  (   (   (   P   P   P            	             �>���   �  @ 	 ;��;�	;uQ;�$;�}Z<��             	                       A�              ?�   �    ?     ?fff?@  ?&ff?    	 @�|g@���@���@�,@�,@�,            C�    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ��~�H?�H��� E�� E��B�           	                                                                                       Ap  ��                      ����BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                    	                                      	     ?��@I�                         	                                      	             ��      Ç               	 C�  D�@ C�                           	 ?��        ?�ؿ��@I�             	 DBTZC5�BjZBa:^B8�@���             	 ��33�ÍC׼��
<#�
?�             	 �H޸��
A�z�BO�V{?�             	 @�ffB233B�B_���L��d�             	 L��J�;�I"�PI?ؒIU߅F�k�             	 L��5K��I��PH�H�I"��F�B             	 L��TK�,kJ��I:�Ie-Gv�l             	                                      	         D�@                          	                                      	         BZ2-                         	         ��                         	         BV-;                         	         ��yR                         	         H��                         	         J��r                         	         J�                         	                                      	         ��                           	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	         ���                         	                                      	         CH                           	         ���                         	         C���                         	         ��;d                         	         @m�                         	         åp�                         	         LΏr                         	         L���                         	         JT�                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 3p$S                    ��������� 	     3b?�                ��������� 	         �@x5            ��������� 	             3�!i        ��������� 	             �7�3��    ��������� 	             � �:�(��3��H��������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	                                      	                                      	                [                     	               e   �                 	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	             �                	            �  c�             	                             	                             	                                 2 E�  E�@     E� D�      Fp         B�  A   A�  C�  D  A   @�                                                                                                      �                                            E�          E�         Fp                                                                                     ?���?ٙ�            	                                
                                                                                                                                                                                                                                                                                          	                   �3��       � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 C`��                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 Cy�f                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      A�XD�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                 ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                             �       F   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$MSKCFMAP  �������                               �$MSKCONREL         �   �$MSKEXCFENB         
�    �$MSKEXCFFNC         
�   �$MSKJOGOVLIM         d�   d�$MSKKEY         �   �$MSKKEY_PANL             �$MSKRUNOVLIM         �   �$MSKSFSPDTYP         
�    �$MSKSIGN         �   �$MSKT1MOTLIM         d�   �$MSK_CE_GRP 1��������  \     	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                             	                                          	                                        �$MSQZ_EDIT      ����    �$MTCOM_CFG 1��������         
       
       
       
       
       
       
       
�$MT_ARC_ENB         �   �$MUAP_CPLENB         �    �$NOCHECK ?�������  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �                  �$NO_WAIT_LN        ���   �$NUM_RSPACE  �������     
   
   
   
   
   
   
   
�$ODRDSP_ENB         �    �$OFFSET_CART         �    �$OFFSET_DIS         �    �$OPEN_FILES     
   ��   
�$OPTION_IO         �   �$OPTM_PRG %�������%$************************************  �$OPWORK ��������    �� �� ��       ���                        	 �                      �      ��$ORG_DSBL  �������                                  �$ORIENTTOL      C�  �A   �$OUT_SIM_DO        �    �$OVRDSLCT ��������    ������   
   
   
   
    �$OVRD_PEXE         �    �$OVRD_RATE         d�   �$OVRD_SETUP ��������     
 ����������������������������������������     
 �����������������������������������������$PARAM2_GRP 1���� 	 d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                                
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                      d                                                                                                                                                                                                                                                                                                                                                                                                                      2                                                                                                                                                                                                          <                                                                                                                                                                                                                                                                                               
                                          P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                  P                                                                                                                                                                                                                                                                                                                                                        	   �  �  �  �  �  �  �  �  �       d 	                                   d 	                                                         	                                                                                                                                                                     �$PARAM_GROUP 1�gX�� `    X, �    �� @D�  D�  ?�  ?�  X,?   ?�      CH  D�  D�                             ;�	l?�   	 ���T��    	 �^� � � � � � � 	 H�kIH��H�+�H���H�{BH&9             	                      	   �  �  �  �  �  �  �  �  � 	 B�  B�  B�  B�  B�  CH                       	 �4    ��Pô  ��  ô               	 �4    ��Pô  ��  ô               	     A6�    ����                 	                      �   �   � 	                                  	   �  �  �  �  F  m  �  �  � 	                                      	  	'� �  �  I� �  ��             	 =���=���=���=���=���=���=���=���=��� 	  @ @ @ @ @ @             	   �  �  �  �  �  �              �    	                                	   ��  ��  ��  ��  ��  ��  ��  ��  �� 	 C4  B�  B�  C�  B�  C�               	 C4  B�  B�  C�  B�  C�                 �C�   	       ���       	        � � I       	 C   C   C   B   B   B                 @   @   @       Dz       	                                      	                                      	                                      	  	'� �  �  I� �  ��            �   � :=             �  @?�ff                                                             	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	  (   (   (   P   P   P            	             �>���   �  @ 	 ;��;�	;uQ;�$;�}Z<��             	                       A�              ?�   �    ?     ?fff?@  ?&ff?    	 @�|g@���@���@�,@�,@�,            C�    ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                       Ap  ��                      ����BH       	                                      	                                      	                                      	 A   A�  A�  A�  A�                      	                                    	                                      	     ?��@I�                         	                                      	             ��      Ç               	 C�  D�@ C�                           	 ?��        ?�ؿ��@I�             	 DBTZC5�BjZBa:^B8�@���             	 ��33�ÍC׼��
<#�
?�             	 �H޸��
A�z�BO�V{?�             	 @�ffB233B�B_���L��d�             	 L��J�;�I"�PI?ؒIU߅F�k�             	 L��5K��I��PH�H�I"��F�B             	 L��TK�,kJ��I:�Ie-Gv�l             	                                      	         D�@                          	                                      	         BZ2-                         	         ��                         	         BV-;                         	         ��yR                         	         H��                         	         J��r                         	         J�                         	                                      	         ��                           	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	         ���                         	                                      	         CH                           	         ���                         	         C���                         	         ��;d                         	         @m�                         	         åp�                         	         LΏr                         	         L���                         	         JT�                          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 3p$S                    ��������� 	     3b?�                ��������� 	         �@x5            ��������� 	             3�!i        ��������� 	             �7�3��    ��������� 	             � �:�(��3��H��������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P         	                                      	 ( 	                                      	                                      	                                      	                                      	                [                     	               e   �                 	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	             �                	            �  c�             	                             	                             	                                 2 E�  E�@     E� D�      Fp         B�  A   A�  C�  D  A   @�                                                                                                                                                                                                                                                                   ?���?ٙ�            	                                
                                                                                                                                                                                                                                                                                          	                   �3��       � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 C`��                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  ��������� 	  � � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 C�                                           	 ��                                   	                                      	                                      	   ,  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	 Cy�f                                 	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J�      � �      � @D�  D�  ?�  ?�   � `?   ?�      C�  D�  D�                             ;�	l?�   	  }�������� 	  } � � � � � � � � 	 F���                                 	                      	   �  �  �  �  �  �  �  �  � 	 D�                                           	                                      	                                      	                                      	    �  �  �  �  �  �  �  �  � 	                             	   �  �  �  �  �  �  �  �  � 	                                      	  +UU                                 	 =���=���=���=���=���=���=���=���=��� 	   ��  �   �   �   �   �   �   �   �  	   &f  &f  &f  &f  &f  &f  &f  &f  &f  �    	                                     	   u0  '  '  '  '  '  '  '  ' 	                                      	                                           ��    	                    	                    	 B                                     @   @   @       ECP      	                                      	                                      	                                      	  +UU                           �     :                ?�                                                               	  �� �� �� �� �� �� �� �� �� 	  8   8   8   8   8   8   8   8   8  >���   �?            	                             	                   �>L��       	 A�                                   	                                       ?�   �    ?�    ?fff?@  ?&ff?    	                                     �     ?�               	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                          ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                                          	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                             	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	                                      	                                                                                                                                	                                      	                                      	                                      	 A   A�  A�  A�  A�                       	                                      	                                    	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������        P 	  P P P P P P P P P          	                                      	 ( 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	 ( 	                             	                             	                             	                             	                             	                             	                             	                             	                                 2                                                                                                                                                                                                                                                                                                                                                        	                                      
                             ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	                   ��{J��$PARAM_MENU ?�������  DEFPULSE              	WAITTMOUT             RCVTMOUT              SHELL_WRK.$CUR_STYLE  SHELL_WRK.$CUR_OPTA   SHELL_WRK.$CUR_OPTB   SHELL_WRK.$CUR_OPTC   SHELL_WRK.$CUR_DECSN  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PASSREL_ID      ���   �    �$PAUSE_PROG %�������%�                                      �$PCCRT         �    �$PCCRT_HOST !�������!PCCRT                             �$PCTP         �    �$PCTP_HOST !�������!PCTP                              �$PC_TIMEOUT      ����   �$PGDEBUG  �������    �$PGINP_FLMSK      ����    �$PGINP_FLTR      ����   �$PGINP_PGATR  �������                     �$PGINP_PGCHK      ����   �$PGINP_TYPE ?������  �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �$PGINP_WORD ?	�������  	FOLGE     	UP        	MAKRO     	SUCHL     	MAKROSP   �$PGTRACECTL 1�������� 
   � �
    � �   � �                                    �$PGTRACEDT Q�������� 
D � 
 5  
 6  
 7  
 8  
 9  
 :  
 ;  
 <  
 =  
 >  
 ?  
 @  
 A  
 B  
 C  
 D  
 E  
 F  
 G  
 H  
 I  
 J  
 K  
 L  
 M  
 N  
 O  
 P  
 Q  
 R  
 S  
 T  
 U  
 V  
 W  
 X  
 Y  
 Z  
 [  
 \  
 ]  
 ^  
 _  
 `  
 a  ��    �   ��    �   �   �   �   �   �   �   �   � 	  � 
  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �    � !  � "  � #  � $  ��    �   �   �   �   �   �   �   �   � 	  � 
  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �    � !  � "  � #  � $  ��    �   ��    �   ��    �   ��    �   ��    �   ��    
 S  
 T  
 U  
 V  
 W  
 X  
 Y  
 Z  
 [  
 \  
 ]  
 ^  
 _  
 `  
 a  ��    
   
   
   
   
   
   
   
   
 	  
 
  
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
    
 !  
 "  
 #  
 $  
 %  
 &  
 '  
 (  
 )  
 *  
 +  
 ,  
 -  
 .  
 /  
 0  
 1  
 2  
 3  
 4   � 

   

   

   

   

   

   

    

 !  

 "  

 #  

 $  

 %  

 &  

 '  

 (  

 )  

 *  

 +  

 ,  

 -  

 .  

 /  

 0  

 1  

 2  

 3  

 4  

 5  

 6  

 7  

 8  

 9  

 :  

 ;  

 <  

 =  

 >  

 ?  

 A  

 B  

 C  

 D  

 E  

 F  

 G  

 H  

 I  

 J  

 K  

 L  

 M  

 N  

 O  

 P  

 Q  

 S  

 T  

 U  

 V  

 W  

 X  

 Y  

 Z  

 [  

 \  

 ]  

 ^  

 _  

 `  

 a  

 b  

 c  

 d  

 e  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  
                            	   
              
 	  
 
  
   ~   ~   
(   
)   
*   
+   
+   
+   
+   
+   
+   �   �   �   �   �   �   �   �   �   �    �   �   �   �   �   

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  

 �  �   � 	  � 
  ~   ~   ~   
   
   
   
   
   
   

   

   

   

   

   

   

   

   

 	  

 
  

   

   

   

   

   

   

   

   

   

   

   

   

   

    �  _   `   a   b   c   d   e   f   g   h   i   j   k   l   m   n   o   p   q   r   s   t   u   v  ��                             	   
                                                                      !   "   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @   A   B   C   D   E   F   G   H   I   J   K   L   M   N   O   P   Q   R   S   T   U   V   W   X   Y   Z   [   \   ]   ^   _   `   a   b   c   d   e   f   g   h   i   j   k   l   m   n   o   p   q   r   s   t   u   v  ��     '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @   A   B   C   D   E   F   G   H   I   J   K   L   M   N   O   P   Q   R   S   T   U   V   W   X   Y   Z   [   \   ]   ^   � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��     � ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    �$PGTRACELEN       ��   ��$PGTRACE_UP ��������   ����$PG_CFG ��������       ����                                                      �$PG_DEFSPD ��������  �     ��$PING_CTRL ��������      8       �$PIPE_CONFIG �����������                   �$PLID_CFG ��������   �$PLID_GRP 1������� �   C�  ��33    B (�H��H�G'4WA�  D	�          �   d      d      d   d   d   d         � 	                                    	                 ´  ´               	                 B�  B�               	                 ´  ´               	                 B�  B�               	                 B
�B�7             	                                      	                 <,1<,1             	                                      	                                      	                                      	                 <,1<,1             	                                      	                                      	                 Dz  Dz                      
 C�q����@�b�?1��                                 	                                      	                                      	                                      	                                      	                 >V̴>WI�             	                                      	                                      	                                        !    
V7.10beta1         @�(�@S33@W�C�    C���C��=B�k�  D�@ D�@ D2ٚ  E��E�D�HC  A�  C  C�  C�  Ap     B�  B�  B�  C�{B&ffB33Bd��B�  B�  BL  B�ffB���BX  �{w�D�An�     ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ���                                                  �   d      d      d   d   d   d          	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                              
                                                  	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                             
V7.10beta1          F@ F@ F@ F@   F@ F@ F@   F@ F@ F@   F@ F@ F@                     ?�     B�  B�                                                               ����$PLID_KNOW_M         �   �$PLID_SV ���������        
                                                                                  	                                      	                                        d      d   d    �$PLIM_GRP 1��������  lC�   	       ���       	        � � I       �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���    	                    	                    �@�    @�  @�  @�    @�  @�  @�    @�  @�  @�    ���$PLMR_GRP 1��������  T        B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�                      B�                   
 B�  B�  B�  B�  B�  B�  B�  B�  B�  B�              �$PLST_GRP1 1�������� 
 0Vacia             Cx:�A+�dA(��A�y�I�H[��IO�Llena             C�q����@�b�?1��            �                  C�                          �                  C�                          �                  C�                          �                  C�                          �                  C�                          �                  C�                          �                  C�                          �                  C�                          �$PLST_GRP2 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP3 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP4 1�������� 
 0�                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �                  �                           �$PLST_GRP5 1��������  0�                  �<                         �$PLST_GRP6 1��������  0�                  �<                         �$PLST_GRP7 1��������  0�                  �<                         �$PLST_GRP8 1��������  0�                  �<                         �$PLST_GRPMAD        �   �$PLST_PARNUM  �������                              �$PLST_SCHMAD         �   
�$PLST_SCHNUM         �   
�$PLST_UPDNUM  �������                          �$PLS_CMP_LIM  ����  '�   �$PLS_ER_CHK  ���� ���    �$PLS_ER_LIM  ����  '�   �$PLS_ER_RST         �    �$PL_MOD         �   �$PL_MOD_ST         �   �$PL_RES_G1 1�������� 
  Cx:�D4f�D4f�C{RHUM
HUM
F�F�   C�qD9�#D9�#Cu�}HY5HY5F�X�                                                                                                                                                                                                                                                           �$PL_RES_G2 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G3 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G4 1�������� 
                                                                                                                                                                                                                                                                                                                        �$PL_RES_G5 1��������                                  �$PL_RES_G6 1��������                                  �$PL_RES_G7 1��������                                  �$PL_RES_G8 1��������                                  �$PL_RES_V 1�������   �  �^�`�^h�]�T�]���$PL_THR_INRT         d�   d�$PL_THR_MASS         d�   Z�$PL_THR_MMNT         d�   Z�$PMON_QUEUE ��������       �      �$PM_GRP 2�������  4      A�  @�                    B�           �$PNS_CUR_LIN        ���    �$PNS_END_CUR         �    �$PNS_END_EXE         �    �$PNS_NUMBER        ���    �$PNS_OPTION         �   �$PNS_PROGRAM %�������%PNS                                   �$PNS_TASK_ID        ���    �$POCFG ��������                                      �$PODATA_GRP 1�������� @ ��   - 2 �����~~����~~�����~~����~~����~~����~~�����~~���~~ 2     " 5     " 5      " 5     " 5     " 5     " 5      " 5    " 5   2                                                    ��    2 ~~���~~�����~~����~~�����~~����~~����~~����~~����� 2     " 5      " 5     " 5      " 5     " 5     " 5     " 5      " 5 2                                                    ��    2 �~~����~~�����~~���~~�����~~����~~�����~~����~~��� 2  5     " 5      " 5    " 5      " 5     " 5      " 5     " 5     " 2                                                    Z    2 ����~~������~~~~������~~����~~������~~����~~����~~ 2    " 5       " 5         " 5     " 5       " 5     " 5     " 5   2                                                   �$POINFO_GRP 1�������� �     �                                                                                                                                                                                                                                                                                                                                                                                                                 �$POIO_GRP 1��������             �$POS_EDIT ��������                               �$POWERFL            �    �$PRGADJ ��������A�  A�  A�  ?   ?   ?      d    �$PRGNS_CFG ��������?�             @   <@�             %�                                                            �$PRGNS_GRP 2�������� �  \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                       \        �   ?�  ?�  A       �t$ �t$ �t$ ****/**/** **:**:**   ****/**/** **:**:**   �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                      �����������������A   �������������                      �                       	                                      	                                      	 �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$ �t$  	                                      	                                     �$PRGNS_PREF ��������      
    �$PRIORITY         ��   ��$PRMPDSPON            �    �$PRMPDSPOUT        �   �    �$PRODUCT_ID �������                       �$PROGGRP_TGL      ����    �$PROTOENT 1��������  (!AF_INET                              !tcp                                  !udp                                  !icmp                                 �$PROXY_CFG ��������  �    )� ****************************************   �)� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** )� **************************************** �$PRO_CFG ��������    %�                                                          ?Lio        ****/**/**/ **:**:**      %�                                         �                        A�    ,  �                                                                                     �$PRO_PREF ��������      
      �$PRPORT_NUM        �   �$PR_CARTREP  �������    �$PSKSTAT         �    �$PSSAVE ��������	2600H621                                              !�                                  !�                                  �                  	�          �        �                         �                      e�                                                                                                      �              !�                                  �$PSSAVE_GRP 1��������     to                  ���������������������$PS_CONFIG ��������                     
          �  �   �v��$PS_CP_CFG 2��������                                                         �$PS_CP_GRP 2�������   �         U�8�?]����㴒Nd���ğ�5�>��?�P�5"D0�|D��D�K    8�?]�����C8���ģ�5�>��?�K�5(D0��D��D�G        8�?�              ?�              ?�                  q8 ��    ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������           ���    ���8����������������������������������������8����������������������������������������    8����������������������������������������       �$PS_MOTION 2�������� 
�                                %�                                      %�                                                                                                                  8�?�              ?�              ?�                                                                                                                                                                                                                                                                                                                             ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �2�%�                                   ��*��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �+z%�                                   �v��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �OO%�                                   &"��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   ��%�                                   �I���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                    ^c%�                                   (�N��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   ���%�                                   +u���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �d�%�                                   >���������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                   �  %�                                   ����������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        ���    ������������%�                                     %�                                     ��������������������������  ������������������  ���������8������������������������������������������������������� ������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������      �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$PURGE_ENBL         �   �$PWFENBDO            �    �$PWF_IO        �   �$PWRUP_DELAY ��������       �$PWR_HOT %������   �%�                                      �$PWR_NORMAL %�������%�                                      �$PWR_SEMI %�������%�                                      �$QSKIP_GRP 1��������  x 	                                      	                                                                              	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ��������������������������������������������������������� 	 ��������������������������� 	 ����������������������������������������������������������$RBTIF      ����    �$RCVTMOUT        ��  ��$RDCR_GRP 1������� � 	 E�*HE�]�    D���D���C�ڜ             	 �t�[��q�)c��5���w�NÊ*             	                                      	 ;��;�	;uQ;�$;�}Z<��                    	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                    	                                      	                                      	                                      	                                             	                                                                                                                                                                                                                                                                                                   �$RDIO_TYPE  �������                                  �$REFPOS1 1�������� 
 x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS2 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS3 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS4 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS5 1��������  x�                                  	                                      	                                         �                                  	                                      	                                         �                                  	                                      	                                         �$REFPOS6 1��������  x�                                  	                                      	                                         �$REFPOS7 1��������  x�                                  	                                      	                                         �$REFPOS8 1��������  x�                                  	                                      	                                         �$REFPOSMASK 1��������     
   
   
   
   
   
   
   
�$REFPOSMAXNO  �������     
                     �$REMOTE  �������   �$REMOTE_CFG ��������          �$REPL_RANGE      ����   �$REPOWER ��������    �$RESM_DRYPRG %�������%�                                      �$RESTART ��������            �$RESUME_PROG %�������%�                                      �$RE_EXEC_ENB         �   �$RGSPD_PREXE         �    �$RGTDB_PREXE         �    �$RGTRM_PREXE         �    �$RMT_MASTER  �������    �$ROBOT_ISOLC  �������                 �$ROBOT_NAME �������KJLTVL111120R01       L T �$ROB_ORD_NUM ?�������  H621  H895 �H895  H895      ���     �             �$RPC_TIMEOUT      ����   x�$RS232_CFG 1��������  LTEACH PENDANT                                  �                  Maintenance Conso                          "   �                  	Unbenutzt                                      �                  	Unbenutzt                                      �                  �$RS232_NPORT        �   �$RSCH_LOG ��������       		RSCH          �$RSMAVAILNUM        ��   �$RSPACE1 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                    ���������  ����������                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE2 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE3 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE4 2�������� 
 �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE5 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE6 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE7 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACE8 2��������  �                                                                                      8�?�              ?�              ?�                                                                                                              �$RSPACEG ��������                           
 
                                                                                  ������������������������������������������������������������                                                                                                              d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������                         d d                                                                                  ������������������������������������������������������������                                             ���������  ���������  ���������  `                  @   @   @                                                                           �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                              �  @   @   @     ���������  ���������  ���������                ����������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  �������������������������������  ���������  ���������  ���������  ��������������������� 
                                         �$RSPACE_MODE  �������    �$RSPACE_S ��������                                                                                                                          	                                     �$RSPCWORK_AD  ��������ܤ�$RSR  �������                  �$RSR_INTVAL        ��    �$RSR_OPTION         �   �$RTCFG ��������                      ?          �  �   �$RV_DATA_GRP 2�������   � D  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  P 	                                      	                                      	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SAF_DO_PULS  ����   �������$SCAN_TIME        ��   �$SCR ����8		      
      
               
                                                                                                                                                                                                                                                                             �         2   2   
   
   d   
   d   2   d                       
 @                                                                          
                               P       
�� @B     T                                                                                    T D��                                                                                                                                                                                                                                                                                                                                                            @                    




                                             @         ;�o             p              
�t� �Di                        �                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                  �                                 0    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                                                                                                                                                                                                  �           �  �  � � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                   T                                                                                                                                                                                                                                                                                                                                                      �                                                       ��                                     	12345678    `!B  �            T                                                                                      T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T BH                                                                                                                                                                                                                                                                                                                                               T :�j                                                                                                                                                                                                                                                                                                                                             T D�                                                                                                                                                                                                                                                                                                                                               T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                  T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   "CH  A�               �          2                   
   d   
  �  	�     2                                                                                                       p  �                                  �                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                                                                                                                                                                                                                                                                                                                                                     �$SCR_GRP 1��� t �            	    � 	    � 	                                  	                                	                                     �      D�@ D�                   �     �                            M-900iA/260L_iC 7890  	M-900iA   	M92C 678      
V06.10         	             
   
   
           	          �       �              	      	          � 	                                                                                                             ��H� 	     	    ��      O����x�@D���D���´  B4�Bp ! 	 Bp ��A���7ej� ´                     =4H��x��D��D��B 	                                                            	                                         	                                     	 B�  B�  BǙ�B�  B�  B�  B�  B�  B�   	 A   A   A   A   A   A   @   @   @    	 @�  @�  @�  @�  @�  @�  ?�  ?�  ?�   	 BH  BH  BH  BH  BH  BH  A   A   A    	 F@ F�` F�`                          	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                            
                                         ?�  @�  @T�                         	 @�  @�  @�  @�  @�  @�  B�  B�  B�  12345678901234567890                                                  A�                	                    	                                                                                                                                           � � � ( ( (                                                        �           	 	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	 B���                                                         	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	 A���                                                         	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �            	          � 	          � 	                                     	                              	 @                                                                      �     �                            Independent Axes 890  		Independe 		Independe     
V06.10         	                              	          �         �               	           	          � 	                                                                                                              ��H� 	     	          ��                                     	                                                              	                                                            	                                          	                                     	 B�  B�  B�  B�  B�  B�  B�  B�  B�   	 @   @   @   @   @   @   @   @   @    	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 A   A   A   A   A   A   A   A   A    	                                      	                                      	                                      	                                      	                                      	                                      	 B�  @   ?�                           	 B�  @   ?�                           	 B�  @   ?�  B�                       	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                             
                                                                              	 @�  B�  B�  B�  B�  B�  B�  B�  B�  12345678901234567890                                                  A�                   	                    	                                                                                                                                                                                                                                �$SEL_DEFAULT        ���   �$SEMIPOWERFL         �   �$SEMIPWFDO         �    �$SERVENT 1�������  L!DUM_EIP                             �j!AF_INET                           !FTP                                  !AF_INET                           !�                                    �!AF_INET                           !RPC_MAIN                            �!AF_INET                           !RPC_VISN                            �!AF_INET                           !TP_INPUT                            �d!AF_INET                           !
PMON_PROXY                          �e!AF_INET                           !TP_PROXY                            �f!AF_INET                           !RDM_SRV                             �g!AF_INET                           !R90                                 �h!AF_INET                           !
RPCM_PROXY                          �i!AF_INET                           !RLSYNC                              8!AF_INET                           !ROSIP                               �4!AF_INET                           !
CETP_MTCOM                          �k!AF_INET                           !	CETP_CONS                           �l!AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           !�                                      !AF_INET                           �$SERVICE_KL ?%������  (%SVCPRG1                               %SVCPRG2                               %SVCPRG3                               %SVCPRG4                               %SVCPRG5                               %SVCPRG6                               %SVCPRG7                               %SVCPRG8                               %SVCPRG9                               %SVCPRG10                              %SVCPRG11                              %SVCPRG12                              %SVCPRG13                              %SVCPRG14                              %SVCPRG15                              %SVCPRG16                              %SVCPRG17                              %SVCPRG18                              %SVCPRG19                              %SVCPRG20                              %SVCPRG21                              %SVCPRG22                              %SVCPRG23                              %SVCPRG24                              %SVCPRG25                              %SVCPRG26                              %SVCPRG27                              %SVCPRG28                              %SVCPRG29                              %SVCPRG30                              �$SERVICE_PRG ?%������  (%                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       %                                       �$SERV_DEV �������MC:           �`��$SERV_MAIL      ����    �$SERV_OUTPUT      ����    �$SERV_REC 1�������   �     	    �   �   �   �   �   �             	                                    	                                	                                     
 �X���6 2     	                    ��������� 	    2    %  �       ��������� 	    T   K����   ~���{���Y��������� 	 �������   G  ����
  ����������X�U'6    	   L  x  N  !  �  ��������� 	       q   �    �   ��������� 	    j����      A�������\��������� 	 ����   �������G���A  ���������X���6      	     s  B  �  �  "���������� 	       A  �      L  ��������� 	 ����   A����   ���������������� 	 ����   ����7���B�����������������XÎ46 2     	    A      Z   L      D��������� 	   �      "      e  ���������� 	 ����   3����   _�������h��������� 	 ����  ����  �����  ����������XÎV6 2     	                      ��������� 	   [   @   2      �  ��������� 	 ����   3����   _�������h��������� 	 ����  �����  ����  	*���������XÎ\6 2     	                     ��������� 	   �   J   2      �  %��������� 	 ����   3����   _�������h��������� 	 ����  }����   �����  	����������X�+�6 2     	    F   $   o   c       X��������� 	   �      %       b  ��������� 	 ����   3����   _�������h��������� 	 ����  ����  ����Q  ����������X�+�6 2     	    '   	      
       ��������� 	   �              �  g��������� 	 ����   3����   _�������h��������� 	 ����  c���7  ����  K���������X�Y�6 2     	                     ��������� 	    4  W    �       #��������� 	    T   K����   ~���{���Y��������� 	 �������   h  j���  %���������X�E�6 2     	                     ��������� 	    ?  ,  �  �       !��������� 	    T   K����   ~���{���Y��������� 	 ��������   �  "����  ����������   	 
 �Vq6 2     	   �    o  �  	q   1��������� 	    1   �  &   -  �    ��������� 	 ����   *�����������I���`��������� 	 ��������   Y  E  �  Y���������W!o6 2     	   <  �  �  �  
   ��������� 	    %   �  H   &  x    ��������� 	 ����   *�����������J���`��������� 	 ������������  G  �  ����������V~u�6 2     	   �  �  Z  �  	9   6��������� 	    0   �  9   8  h    ��������� 	 ����   *�����������I���`��������� 	 �������3   ,  �  �  ����������VvC6 2     	   =  �  �  �  
   ��������� 	    (   �  K   *  �    ��������� 	 ����   *�����������J���`��������� 	 ���)��������  B  �  Q���������U�Mc6 2     	   /  j  �  �  	�   !��������� 	    /   �  x     V    ��������� 	 ����   *�����������J���`��������� 	 ������������  )  �  e���������W��86 2     	   k  �  �  �  
5   ��������� 	       �  K   *  �    ��������� 	 ����   *�����������J���`��������� 	 ���A���9���_  �  d  7���������W~`V6 2     	   ,  p  �  �  	�    ��������� 	    ,   �  4   +  �    ��������� 	 ����   *�����������J���`��������� 	 ����������t  �  �  !���������W}`6 2     	     Y  �  �  	�   %��������� 	    *   �  4   6  �    ��������� 	 ����   *�����������J���`��������� 	 ���t��������  �  c  ����������X#-#6 2     	     X  �  �  	�   %��������� 	       �  3   9  �    ��������� 	 ����   *�����������J���`��������� 	 ������������  ]  +  ����������L|��6 2    	       
      *   U    ��������� 	   =   �    �   :  x��������� 	 ����   0����   V�������`��������� 	 ���y  ���  z���i  Q���������   s 	                                     	                                      	                                     	                                      
 �W}l46 2     	   ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������W�M�6 2     	   p������������������������ 	     ������������������������ 	   (������������������������� 	     ������������������������X#-#6 2     	   ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������X,D�6 2     	   ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������XJ��6    	   "i������������������������ 	     ������������������������ 	   P������������������������� 	     ������������������������V�(�6 2     	   D������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������V�86 2     	   ;������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������W!o6 2     	   k������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������WT��6 2     	   ^������������������������ 	     ������������������������ 	   (������������������������� 	     ������������������������Wa1�6 2     	   ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������    
 �Vq6 2     	   	M������������������������ 	     ������������������������ 	   (������������������������� 	     ������������������������W!o6 2     	   k������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������V~u�6 2     	   p������������������������ 	     ������������������������ 	   (������������������������� 	     ������������������������VvC6 2     	   y������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������U�Mc6 2     	   9������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������W��86 2     	   ������������������������� 	     ������������������������ 	   (X������������������������ 	     ������������������������W}`6 2     	    ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������L|��6 2    	     ������������������������ 	     ������������������������ 	   ������������������������� 	     ������������������������X#-#6 2     	   ������������������������� 	     ������������������������ 	   (������������������������� 	     ������������������������V��6 2     	   #W������������������������ 	     ������������������������ 	   (������������������������� 	     ������������������������   � 	                                     	                                      	                                      	                                      
 �U&�v6 2     	   ������������������������� 	     ������������������������ 	   ������������������������� 	     ������������������������UZK<6 2     	   ������������������������� 	     ������������������������ 	   ������������������������ 	     ��������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������    
 �Vq6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������W!o6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������V~u�6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������VvC6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������U�Mc6 2     	   ������������������������� 	     ������������������������ 	   '������������������������ 	     ������������������������W��86 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������W}`6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������L|��6 2    	     ������������������������ 	     ������������������������ 	   '������������������������� 	     ������������������������X#-#6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������V��6 2     	     ������������������������ 	     ������������������������ 	   '������������������������ 	     ������������������������     	                                      	                                      	                                      	                                      
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������     
 ���������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_RV 1�������   �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ����������������������������$SERV_TOP10 1�������   � 
 6 2   �6    a6�   6    6 *   6�   6    C6�   6r _   6 s   �$SERV_TYPE      ����    �$SHELL_CFG ��������                                                                %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                   %RSR                                                       �  �   %                                                                                                     �         �   2   d                                �$SHELL_CHK 1��������                                                                                                                                                                                                                                                                                                                                                                                  �$SHELL_COMM ��������                        �$SHFTOV_ENB         �    �$SHOW_REG_UI         �    �$SIMWAITENB            �    �$SIMWAITOUT        �   �    �$SIMWAITTIM       ��   �    �$SIMWAITVAL            �    �$SI_UNIT_ENB         �   �$SLC_RETRY         �   �$SMB_HDDN 2��������    ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  ������������������������  �������������������������$SMON_ALIAS ?e������ ( he�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      e�                                                                                                      �$SMON_DEFPRO ������ *SYSTEM*    ��$SMON_RECALL ?}������ ( �}�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              }�                                                                                                                              �$SNPX_ASG 1�������� P 0 '%R[1]@1.1                              ?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    � ?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    � ?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    � ?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    � ?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    ��?�      %                                    9v ?�      %                                      ?�  �$SNPX_PARAM ��������  �	�             P                           ��$SOFT_KB_CFG        ���    �$SOPIN_SIM  �������                                                  �$SRVQSTP_DSB  �������                                  �$SSR ������� � & FOLGE011 .......................0046        �$STHI_CHANGE         �    �$STHI_GRPNUM         �    �$STOP_ON_ERR         �    �$STOP_PTN ������C �$STRING_PRM         �   �$SVDT_GRP 1�������    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                    	                   �$SVPRG_COUNT        ��    �$SVPRG_ENB         �    �$SVPRM_ENB         �    �$SVPRM_UPD 1������� T  
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                      
                     �$SV_CTRL_NUM        
�   �$SV_GUN_CTRL 2��������                 /   /   
               4   4   
                        
                           
                           
�$SYSDEBUG  ����   d�    �$SYSDSP_PASS       B?�    �$SYSLOG ��������         �^��                      �       UD1:\SYSLOG               �$SYSLOG_MPC ��������                                    �       UD1:\SYSLOG2              �$SYSLOG_SAV ��������                     UD1:\SYSLOGSV         �$SYSTEM_TIME 1��������  ( @�     0��        �e                 @�     0��        �O                 @�     0��        �O                 @�     0��        �H                �$T1SVGUNSPD        '�   ��$TASK_OPTION  ������   �   �$TA_DISP_ENB         �    �$TBCCFG ��������                                                 `                             	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                                                                	                                      	                                      	                                         ��������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������������  ���������  ���������  ��������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������    �$TBCSG_GRP 2��������  �     
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   
 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ��� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ��������������������������������� 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������ 
 ������������������������������A��*SYSTEM*   V8.2306       4/24/2014 A t  *SYSTEM* *SYSTEM*  F�TBCPARAM_T   �$MC_MAX_TRQ  $MAX_TRQ_MGN  $MC_GRAV_MGN  $MC_STAL_MGN  $MC_BRK_MGN  $MC_NOLD_MGN  $SHORTMO_LIM  $SHORTMO_MGN  $MC_NOLD_TRQ  $J_LIN  $SPL1  $SPL2  $SPL3  $SPL4  $SPL5  $SPL6  $SPL7  $SPL8   ��TBC_GRP_T � $TBC_ACCEL1  $TBC_ACCEL2  $TBC_PATH1  $TBC_PATH2  $PATH_RATIO  $TBC_PARAM 2  	$CNT_SCALE  $SHORTMO_SCL  $MIN_ACC_UCA  $MIN_CAT_UMA  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2L_UPR_ANG  $J2L_LWR_ANG  $J2L_UPR_MGN  $J2L_LWR_MGN  $R_F2LSHRT  $R_F2LLONG  $MIN_F2LSHRT  $MIN_F2LLONG  $MIN_ACRL_S  $MIN_ACRL_L  $MIN_PAYLOAD  $HVAL   $HMGN   $FLEXL   ��TBJ_ACC_T  :$ACC_LEN1  $ACC_LEN2  $DEC_LEN1  $DEC_LEN2  $ACCEL_RATIO  $DECEL_RATIO  $SLOW_AXIS  $F1ACC_I  $F2ACC_I  $F1DEC_I  $F2DEC_I  $MOVE_TIME  $S_INERTIA   	$D_INERTIA   	$TORQUE_ACC   	$TORQUE_DEC   	$DISPLACEMNT   	$ACCTIME   	$DECTIME   	$VEL_MAX_ACC   	$VEL_MAX_DEC   	$VEL_TCV_ACC   	$VEL_TCV_DEC   	$TRQ_TCV_ACC   	$TRQ_TCV_DEC   	$TRQSTAT_ACC   	$TRQSTAT_DEC   	$J_STAT_ACC   	$J_STAT_DEC   	$M_STAT_ACC  $M_STAT_DEC  $J_MODE  $DT_ACC   $DT_DEC   $ACC2_STP   $DEC2_STP   $AT_MODE  $AT_AXS   	$AC_ACC   	$AC_DEC   	$JK_ACC   	$JK_DEC   	$VK1  $VK2  $VK3  $JJ0  $JJ1  $JJ2  $JJ3  $AA1  $AA2  $AA3  $AA4  $AA5  $TRQ_N1_ACC   	$TRQ_N1_DEC   	$VEL_MAX   	$LINE_NUM  l�TBJCFG_T  � $GROUP_MASK  $MB_CONFLICT  $MB_REQUIRED  $DEBUG  $UPDATE_TIME  $TBJ_SELECT  $TBJ_STAT   $TJ 2 $JERK_CTRL  $MOTN_INF  $TBJ_DEBUG  $HAND_VB   �TBJOP_GRP_T  $ $F2MGN  $MINF2  $COMP_SW   ��TBPARAM_T � $$MR_MAX_TRQ  $MR_STAL_TRQ  $MR_BRK_TRQ  $MR_BRK_VEL  $MR_NOLD_VEL  $MA_LOAD_TRQ  $MD_LOAD_TRQ  $MAX_TRQ_MGN  $MA_GRAV_MGN  $MA_STAL_MGN  $MA_BRK_MGN  $MA_NOLD_MGN  $MD_GRAV_MGN  $MD_STAL_MGN  $MD_BRK_MGN  $MD_NOLD_MGN  $PTH_GRV_MGN  $PTH_STL_MGN  $PTH_BRK_MGN  $PTH_NLD_MGN  $DYN_FRC_MGN  $MR_NOLD_TRQ  $R_ACC_MGN  $R_DEC_MGN  $R_LONG_MGN  $J_ACC  $J_DEC  $DT_MGN  $SP1  $SP2  $SP3  $SP4  $SP5  $SP6  $SP7  $SP8  T��TBJ_GRP_T   $$TBJ_ACCEL1   	$TBJ_ACCEL2   	$ASYM_PARAM   $TB_PARAM 2 	$SHORTMO_SCL  $LONGMO_SCL  $MIN_ACC_SHM  $MIN_ACC_UMA  $SHORTMO_MGN  $LONGMO_MGN  $MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	$PAYLOAD_MGN  $J2J_UPR_ANG  $J2J_LWR_ANG  $J2J_UPR_MGN  $J2J_LWR_MGN  $INERTIA_VIB   $INERTIA_VI2   $IV_UNIT  $IV_UNIT2  $R_F2JACC  $R_F2JDEC  $R_F2JLONG  $MIN_F2JACC  $MIN_F2JDEC  $MIN_F2JLONG  $MIN_ACRJ_S  $MIN_ACRJ_L  $MIN_PAYLOAD  $HVAL   $HMGN   $HAXS   $FLEX    ��TCPPIR_T    $ENABLE_TCPP  $TCDELAY    ��TCPPSPEED_T  X $TCDELAY_MON  $VSPEED  $SPEED  $ACCEL  $TIMESTAMP  $PROG_SPEED  $MOTYPE  �TCPP_CFG_T 	 | $NUM_TCPPSEG  $GROUP_NUM  $TCPP_TIME  $WARNING_ENB  $OTF_TIM_ENB  $DEBUG_TASK  $DEBUG_MAIN  $TCPP_CMP_SW  ��TCPSPDCFG_T 
 � $TCDELAY  $HEARTBEAT  $SETUP_CFG  $SPD_MARGIN  $DEBUGFLG1  $DEBUGFLG2  $SPARE_STR1 $SPARE_STR2 $SPARE_LONG1  $SPARE_LONG2  $SPARE_REAL1  $SPARE_REAL2  ��TCPSPDOUT_T  p $ENABLE  $TARGET_TYPE  $TARGET_IDX  $MIN_VALUE  $MAX_VALUE  $MIN_SPEED  $MAX_SPEED  $GROUP_NO  �TP_THR_TABLE  $ $THR_ENB  $DI_NO  $DO_NO   ��THR_CFG_T  0 $MAX_IO_SCAN  $MIN_SCAN_TI  $SCAN_TIME  ��TIMER_T  � $COMMENT $TIMER_VAL  $STR_EPT_IDX  $STR_LIN_NUM  $END_EPT_IDX  $END_LIN_NUM  $TID_NUM  $DUMMY13  $PS_OVERFLOW   $OVERFLOW  $FLAG_TYPE  $FLAG_IDX  $GLB_TMR_ENB  $GLB_TMR_STR  ��TORQCTRL_T  X $DEBUG  $GRP_STT   $SBR_PAM21_V   T$SV_ERR_MOD   $SV_ERR_CLR   $ACTION  �TPGL_VIEW_T  4 $X  $Y  $Z  $WZ  $P  $R  $CAMERA    ��TPGL_UVIEW_T   $NAME $GIF }$VIEW �TPGL_CAM_T  L $NAME $ID }$FID E$GIF }$NEARPLANE  $FARPLANE  $DISTANCE    ��JOG_RAD_T   $JOINTS   	 �TPGL_MSET_T    $NAME E$ID }$TIMECONST  8�TPGL_CONF_T � $MOUNT ?� $LOCK_FOLLOW  $DBGLVL  $GLDBGLVL  $TEST_XML }$TEMPINT   $TEMPSTR ?� $USER_VIEWS 2 $CAMERAS 2 $TEMP_LOCS 2 $SCENE_VIEW 2  $KAREL_TMO  $TPDRAW_TMO  $JOG_VECLEN  $JOG_RADIUS 2 $CHECK_TOOLS  $CHECK_VIS  $REG_VIS32  $REG_VIS64  $MACHSET 2 $CONT_IDX  $DUMMY29  $VISIBLE   @$RAIL_BOXES   $ROBOT_XML ?� $SHOWWARN   $PS_CONTROLM   $CONTROLMAX  $CONTROLMASK   $FP_TO_FK ! U��TPGLMACH_T   $JOINTS   	`�RECLOC_T   $SLOTS !  ��TPGL_OUT_T  X $VIEWS 2 $SELECTED ?� $PIP_XML }$NODEVIS   @$MACHINES 2 $RECORDEDLOC 2 �TPP_MON_T  D $GLOBAL_MT  $LOCAL_MT  $MON_NUM  $GMON_TID  $SYSMON_ADR  �TPSTRTCHK_T  , $ENABLE  $ALLOW_NAME $ALLOW_LINE   ��TPVWVAR_T  � $TPVIEW_ENB  $PREV_RTN  $EDIT_RTN  $VSHWRK  $DEBUG  $DISPLAY  $INDENT1  $INDENT2  $HEAD1 $HEAD2 $EDIT_KEY  $TCPSPD_KEY  $JMPCALL_ENB  d�TRACE_CFG_T  D $ENABLE  $ITEMS  $CHANNELS  $DEBUG  $TICKS  $MIN_MM  ��TRACE_CHNL_T  @ $ITEM_NUM  $TCP_GP_NUM  $VISIBLE  $STYLE  $COLOR   �TRACE_ITEM_T  t 
$PRG_NAME %$VAR_NAME =$DESC !$UNITS $TYPE  $IO_TYPE  $PORT_NUM  $SQUARE  $SLOPE  $INTERCEPT  '�TSCFG_T  $GRP_MASK  $MODE_MASK  $STATUS  $OPT_VAL  $SIZE  $FNAME_TYPE  $PS_PROC   $PROC  $OUTPUT  $OUTPUT_DONE  $AXS_MSK_ENB  $AXIS_MASK   $CUR_RECTIME  $TOT_CHN_NUM  $MINFREQ_US  $SETFREQ_POW  $LPARAM   
$FPARAM   
$PATH_NAM $DUMMY19  $DUMMY20   l�TSR_GRP_T  l $MR_MAX_TRQ   	$MR_STAL_TRQ   	$MR_BRK_TRQ   	$MR_BRK_VEL   	$MR_NOLD_VEL   	$MA_LOAD_TRQ   	$MD_LOAD_TRQ   	$MA_GRAV_MGN   	$MA_STAL_MGN   	$MA_BRK_MGN   	$MD_GRAV_MGN   	$MD_STAL_MGN   	$MD_BRK_MGN   	$MJ_ACC_MGN   	$MC_ACC_MGN   	$MC_STAL_MGN   	$MC_BRK_MGN   	$MIN_CYC_ID 	$MIN_C_ID_E1 	$MIN_C_ID_E2 	$MIN_C_ID_E3 	�TSSCB_T ! h $DSP_NO  $DSPAX_NO  $DATA_SEL  $OUT_CHANNEL  $ADDRESS  $BIT_SHIFT  $USE_2CH  $MONITOR  �TXSCREEN_T " $ $DESTINATION }$SCREEN_NAME  L�REQ_DATA_T # T $ERR_TYPE  $ERR_GRP  $ERR_AXIS  $AXIS_TYPE  $ERROR_DIST  $ERR_TIME    �UECFG_T $ � 	$CHK_VERSION  $RSM_CHK_ENB  $UNEXCEP_ENB  $RSM_THRS_R  $RSM_THRS_L  $UNEX_THRS_R  $UNEX_THRS_L  $REQ_COUNT  $REQ_DATA 1# 
�UEGRP_T % 0 $ERR_COUNT  $PROGMTN_FLG  $CURR_POS   	��UI_MENHIS_T & 8 $HIST_HEAD  $HIST_ENTRY ?� $DUMMY2  $DUMMY3  �UI_MOUSE_T ' @ $ACTION  $BUTTON  $ROW  $COLUMN  $TIME  $RESERVED  �UI_PANEDAT_T ( � $PAGEURL }$FRAME )$HELPURL }$PARAMETER1 )$PARAMETER2 )$PARAMETER3 )$PARAMETER4 )$PARAMETER5 )$PARAMETER6 )$PARAMETER7 )$PARAMETER8 )$INTERVAL  $PANESTATE  $DUMMY14  $MOUSE '�UI_USRVIEW_T ) < $MENU $CONFIG $FOCUS $PRIM m$DUAL m$TRIPLE m�UNDO_CFG_T *  $UNDO_ENB  $WARN_ENB  L�USER_INFO_T + 8 $USR_PROG %$TASK_ID  $USR_POSIDX  $USR_PR_USE  �USER_TOOL_T , 4 $X  $Y  $Z  $W  $P  $R  $TOOL_NUM  }�USER_UFRAM_T - 4 $X  $Y  $Z  $W  $P  $R  $UFRAME_NUM  �USER_OFFST_T . D $TOOL_OFST 1, $UFRAME_OFST 1- $GUN_WIDTH   $ENB_SUBNUM   
�USRTOL_GRP_T / @ $DIST_TOL  $ORNT_TOL  $RAUX_TOL  $TAUX_TOL  $ENABLE  �VCCM_CFG_T 0  $SC36MFB1ENB  ���VCMR_CAM_T 1h $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DETECT_TYPE  $DRIVE_TYPE  $SET_VTCP  $DEBUG_CODE  $DMY_UBYTE  $CAMERA_NAME %$DISTORTION1  $DISTORTION2  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $HANDEYE  $EXPOS_TIME  $NUM_MUL_EXP  $FOCAL_DIST  $GD_SPACING  $TRGT_DIST  $TRGT_W  $TRGT_P  $TRGT_R  $NUM_RETRY  $UTOOL   ��VCMR_TRGT_T 2  $TARGET_PNT   	t�VCMR_CRPR_T 3 d $AXIS_FLAG   	$NUM_AXS_REP  $SWING_ANG   $NUM_MS_POSE  $BASE_POSE   	$EVALUE_IDX   ��VCMR_CHKM_T 4 @ $EVALUE_IDX  $MAX_MS_ERR  $MEAN_MS_ERR  $WORST_POSE   ��VCMR_MRCV_T 5 � $ORG_MST_CT   	$ORG_UFRAME   $ORG_REF_POS   	$ORG_REF_CT   	$RCV_ANG_PAM   	$NEW_MST_CT   	$NEW_UFRAME   $NEW_REF_POS   	$NEW_REF_CT   	$EVALUE_IDX  $MAX_RC_ERR  $MEAN_RC_ERR  $WORST_POSE  $MASTER_TIME  $DEBUG_MODE   ��VCMR_GRP_T 6 � $STAT_FLAGS  $MENU_CODE  $GROUP_NUM  $UTOOL_NUM  $CAMERA 1$TARGET_ID 22 $CREATE_PRG 3$DATA_ID  $CHK_RESULT 4$RECOVERY 5$EXT_INT1  $EXT_INT2  $EXT_INT3  $EXT_INT4  $EXT_REAL1  $EXT_REAL2  $EXT_REAL3  $EXT_REAL4  �VISION_CFG_T 70 &$DATA_PATH  $DATA_CACHE  $LOG_PATH  $LOG_EXPATH  $LOG_TIMEOUT  $MC_LIMIT  $FR_LIMIT  $TD_LIMIT  $DEBUG_MODE  $HOST_NAME  $COMM_PORT  $ROBOT_NAME  $FLAGS  $MAX_PAGES  $MIN_VPOOL  $VPOOL_SZ32  $VPOOL_SZ64  $VPOOL_SZ128  $VPOOL_SZCAL  $VPOOL_LIM  $VPOOL_WAIT  $TMPPOOL_LIM  $FAILIMG_IDX  $LOADIMG_IDX  $NUM_IMREGS  $IMREG_SIZE  $GPM_CANDMAX  $NUM_ASYNBUF  $NUM_VRTDBUF  $VRTDBUF_SIZ  $TOLE_2D_Z  $TOLE_2D_WP  $PC_SETUP  $LOGQUE_MAX  $ECCU_RETRY  $VEMT_PATH  $VEMT_LIMIT  $VIRCIMG_SIZ  �VISION_GRP_T 8  $BACKLASH   	�VLEXE_CFG_T 9 D $ENABLED  $DATE  $FLDR_INDEX  $FILE_INDEX  $REC_INDEX  �t�CUSTOMMENU_T : $ $TITLE $PROG_NAME %$OPTION  �VSHIFT_CFG_T ;` $DATA_NAME 	$CAMERA_NAME %$EXPOSURE  $WIN_RADIUS  $WIN_POS_X  $WIN_POS_Y  $DISP_SCALE  $DISP_LUT  $OUTPUT_BMP  $LIM_DIST  $LIM_ANGLE  $LIM_TILT  $LIM_SCORE  $LIM_CNTRST  $WARN_DIST  $WARN_ANGLE  $WARN_TILT  $WARN_SCORE  $WARN_CNTRST  $VISION_TYPE  $CAMERA_TYPE  $CAMERA_PORT  $DUMMY23  $USED_CAMTYP   l�VSMO_CFG_T <  $ENABLE  $ADJUST_TIME  �WAIT_DATA_T =  $PROG_NAME %$LINE_NUM  �WV_AXSRST_T >   $AXIS_MASK  $THRESHOLD   %�ZABC_GRP_T ?  $ZABC_MODE   
 p�ZMPCF_GRP_T @   $ZMP_ENB  $ZMP_DMY_LNK   
��ZMPOS_GRP_T A � $M_POS_ENB  $CMCMD_SCL  $CART_MCMD   	$P_ACT $J_ACT   	$P_DES $J_DES   	$P_DES2 $J_DES2   	$UXWPR_ENB  $UXEUL_ENB  $UXWPR_ACT   $UXWPR_DES   $UXEUL_ACT   $UXEUL_DES    ���ZP_CFG_T B  $ENABLE  $DEBUG  P�ZP_CYLINDER_ C 8 $RADIUS  $HEIGHT  $PROG_NAME ?( $LINE_NUM   2��ZP_GRP_T D � $OPTIONS   
$BREAK_TIME  $WORK_SHIFT  $ENABLE  $RV_LIFE   	$SHIFT_OVC   	$PART_ID  $OPTM_RATE   
$MAX_I_RATE  $MAX_DI_RATE  $TRACE_ENV  t�ZP_SPHERE_T E , $RADIUS  $PROG_NAME ?( $LINE_NUM   l�$TBC_GRP 2������� dX,X,?    	 HD|� ?�  ?�  ?L��?L��?L��?�  ?�  D� A                                   D�@ ?�  ?�  ?L��?L��?L��?�  ?�  D  BH                                  D�@ ?�  ?�  ?L��?L��?L��?�  ?�  D  B                                   C  ?�  ?�  ?fff?fff?fff?�  ?�  CB  B�                                  C  ?�  ?�  ?L��?L��?L��?�  ?�  CB  Bp                                  C  ?�  ?�  ?fff?fff?fff?�  ?�  CB  B�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  @   ?�  ?�  ?�  ?�      ?�  ?�      ?�                                  ?L��?�     P   P	V3.00     	m92c      	****      	�          BH                  ?�ff?���   x   d?�  ?�                                            ?�  BH                                          ������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  ������������������������������������������� 	 H������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ������������������������������������  ������������  ������������  �������������������������������������$TBJCFG �������                 �                                     �                                                 	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                      	                                                                                                              	                                      	                                      	                                      	                                      	                                                                                      	                                      	                                      	                                         ������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������������������������������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������������  ���������  ���������  ���������  ������������ 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������������������������������������������� 	 ��������������������������� 	 ��������������������������� 	 ������������������������������                                             �$TBJOP_GRP 2�������  ?���Cz     	����������������������������$TBJ_GRP 2������� � 	  �X�X�       	 �^, �,�        @   ?�   	 �D|� D|� D|� CQffC�s3        ?�  ?�  ?��?��?   ?�  ?��?��?   ?�  ?L��?L��?L��<SZ�D�3@   @�  @   B4  A�      ?�                              D�� D�� D�� C�C�s3        ?�  ?�  ?L��?L��?L��?�  ?L��?L��?L��?�  ?L��?L��?L��;�t�D�?�  @   ?�  B�  A�      ?�                              D�� D�� D�� C�C�s3        ?�  ?�  ?L��?L��?L��?�  ?L��?L��?L��?�  ?L��?L��?L��;�t�D�?333?�  ?fffB�  B       ?�                              C�C�C�C���C�s3        ?�  ?�  ?333?333?   ?�  ?333?333?   ?�  ?333?333?   ;���CA�f?&ff?@  ?�  CR  B�                                      C�C�C�C���C�s3        ?�  ?�  ?L��?L��?��?�  ?L��?L��?��?�  ?L��?L��?��;�8CA�f?fff?���?���B�  Bp                                      C�C�C�C���C�s3        ?�  ?�  ?fff?fff?��?�  ?fff?fff?��?�  ?fff?fff?��=%CA�f?��?�  ?�  C>  B�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      ?�  ?�  ?�  ?�  ?�          ?�  ?�  ?�  ?�      ?�  ?�  ?�      ?�  ?�  ?�              ?�  ?�  ?�  ?�  ?�                                      C�         P   P?�  ?�  	V3.00     	m92c      	****      	�          BH                    F� G G'& GA2 G[= GuH G�� G���G���G�� G���G�ƀG�/ HX�H+ HA�@HX��Ho]�H��H�p                                   C�� Gk G�h�H/�@Hj H�@`H�w�H̯@H��I� I*�I �p=���<���?�  ?�  ?�     n   �   (?�  ?�                                                          ?���@   ?�  ?�                               	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  ������������������������������������ 	 ��������� 	 ���������  ������ 	 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������	�          	�          	�          	�          ���������������  ������������������������������������������������������������  ���������������������������������������������������������������������������������������������  ������������  ������������  ����  �������������������������������������$TCPPACTSW  ������    �$TCPPIR �������   CH  �$TCPPSPEED ������ CH                      UD�     �$TCPP_CFG 	�������                          �$TCP_SPD_CFG 
�������      	�   :�o        �              �                              �$TCP_SPD_NUM      ����   
�$TCP_SPD_OUT 2������� 
                                                                                                                                                                                                                                                                                                              �$TCZEROSPD              �$TESTPARS  ������   �    �$THRESTABLE 1�������                                                                                                 	           
                                                                      �$THRRDITABLE 1�������                                                                                          �$THRRDOTABLE 1�������                                                                                          �$THRSDITABLE 1�������                                                                                                                                                                                                                                                                                                                                                                                                   �$THRSITABLE 1�������                                                                                                             	           
                                                           �$THRTABLENUM  �������          �$THR_CFG �������   
   @   `�$TIMEBF_TTS         
�   �$TIMEBF_VER        
�   �$TIMER 1�������   8�                    �4 ��  H��         �      �                   � �  ��         �       �                    �0� 
Z  ��         �       �                     � 
  ��         �       �                    C�� 
+  ��         �       �                    �� �  ��         �       �                   �g���  H��         �      �                   �g���  H��         �      �                   <g ��  H��         �      �                    
T ��  H��         �      �               ��w    g�g� ��         �       �               �oX    �  �   ��         �       �               �CP    �  �   ��         �       �               Y    �  �   ��         �       �               �Ϫ    �  �   ��         �       �               ?fN    �  �   ��         �       �               ��l    �  �   ��         �       �               ��I    �  �   ��         �       �               ?�    �  �   ��         �       �               ��    �  �   ��                   �               ��    �  �   ��                   �               UTO    �  �   ��                   �                      �  �   ��                   �                      �  �   ��                   �               �     �  �   ��                   �                I    �  �   ��                   �                   �  �   ��                   �                      �  �   ��                   �                      �  �   ��                   �                �    �  �   ��                   �                    �  �   ��                   �                      �  �   ��                   �$TIMER_NUM        @�    �$TMI_CHAN          �    �$TMI_DBGLVL         �    �$TMI_ETHERAD ?�������  0000:e0:e4:34:13:7f 0000:e0:e4:34:13:80 �                  0000:e0:e4:34:13:82 �$TMI_ROUTER !�������!ROUTER                            �$TMI_SNMASK ?�������  255.255.255.0     255.255.255.0     255.255.255.0     255.255.255.0     �$TOOLOFS_DIS         �    �$TORQCTRL ������                                       T                                                                                                                                                                                                                                                                                                                                                                                                                         �$TPE_DETAIL         �   �$TPGL_CONFIG ������  �?/cell/$CID$/grp1              ?�                                                                                                  �/cell/$CID$/grp2                                                                                                                  �/cell/$CID$/grp3                                                                                                                  �/cell/$CID$/grp4                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                             }�                                                                                                                                                                                  ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                    �User View 1           }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345 ���������������������User View 2           }�                                                                                                                              ���������������������User View 3           }�                                                                                                                              ���������������������User View 4           }�                                                                                                                              ���������������������User View 5           }�                                                                                                                              ���������������������User View 6           }�                                                                                                                              ���������������������User View 7           }�                                                                                                                              ���������������������User View 8           }�                                                                                                                              ��������������������� lCamera 1              }�                                                                                                                              E�                                                                      }}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345             Camera 2              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 3              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 4              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 5              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 6              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 7              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 8              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������Camera 9              }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 10             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 11             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 12             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 13             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 14             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 15             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������	Camera 16             }�                                                                                                                              E�                                                                      }�                                                                                                                              ���������  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������                               ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   
   (  �  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������                 �E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ���E�                                                                      }�                                                                                                                              ����� @ ����������������������������������������������������������������  ��������  ��*frh:\tpgl\robots\m900ia\m900ia_260l_ic.xml                                                                                                                                                                                                                � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          � frh:\tpgl\robots\dummy\dummy.xml                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                          ��                                                                                                                                                                                                                                                            ���������     ����������������  88�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  8�?�              ?�              ?�                  �$TPGL_OUTPUT ������   ���?�              ?�              ?�                  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ��  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �  2345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     �}12345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345     }�                                                                                                                               @ ����������������������������������������������������������������  ( 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ��������������������������� 	 ���������������������������  �  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8����������������������������������������  88����������������������������������������8����������������������������������������8�����������������������������������������$TPOFF_LIM      ����   �$TPON_SVOFF         �    �$TPP_MON �������          2        �$TPSTRTCHK �������    �                  �$TPVTCOMPAT         �    �$TPVWVAR �������                   �                  �                       �$TP_DEFPROG %�������%FOLGE011                              �$TP_DISPLAY  �������    �$TP_INST_MSK  �������          �$TP_INUSER         �    �$TP_LCKUSER         �    �$TP_QUICKMEN         �    �$TP_SCREEN �������tpsc  �$TP_USERSCRN �������t_sc  �$TP_USESTAT         �    �$TRACE_CFG ������         	       
?�  �$TRACE_CHNL 2������ 	                 �                 �                 �                 �                 �                 �                 �                 �                 � �$TRACE_ITEM 2������  �%$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          %$123456789012345678901234567890123456  =<123456789012345678901234567890123456789012345678901234567890  !123456789012345678901234567890    1234567890123456                          �$TSCFG ������                 �  �                                                   
                                          
                                         UD1:\               ���$TSR_GRP 1 ������ � 	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678   	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @   @   @   @   @   @   @   @   @    	 @�  @�  @�  @�  @�  @�  @�  @�  @�   	                                      	                                      	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�   	 ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  	12345678  	12345678  	12345678  	12345678  �$TSSCB 2!������                                                                                                                                                                                                  �$TX_SCREEN 1"������ 
 �}ipnl/pnlgen.htm                                                                                                               Panel setup               }	index.STM                                                                                                                     
Robot Info e              }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          }�                                                                                                                              �                          �$UALRM_MSG ?������� 
  �                              �                              �                              �                              �                              �                              �                              �                              �                              �                              �$UALRM_SEV  ������� 
   �$UECFG $������           @�  A�  A   B�   QW 
   �         A B�X�u  �         A =8X  �         A >�X��  �         A >eX��  �         A <EX�  �         A C�X  �         A EcX��  �         A EX�  �         A BX�+  �         A A�X�P�$UEGRP 2%������  0 Q     	 ?�
��
�?
�4�2���9���                    	 B�                                    %     	 B�                                          	                                     �$UI_DEFPROG ?%�������  (%MAKRO050 .......................0002  %MOTN005  .......................0001  %�                                      %�                                      %�                                      %�                                      %�                                      %�                                      �$UI_INUSER  �������                                  �$UI_MENHIST 1&������  (   ��-/SOFTPART/GENLINK?current=editpage,MAKRO050,1                                                                                     �'/SOFTPART/GENLINK?current=menupage,37,1 011,40                                                                                    �(/SOFTPART/GENLINK?current=menupage,381,1 25,1 .....................0019,1                                                         �(/SOFTPART/GENLINK?current=menupage,190,1 20,90                                                                                    �(/SOFTPART/GENLINK?current=menupage,153,1 25,1                                                                                     �-/SOFTPART/GENLINK?current=editpage,FOLGE125,5                                                                                     �-/SOFTPART/GENLINK?current=editpage,FOLGE011,1                                                                                     �'/SOFTPART/GENLINK?current=menupage,23,1  25,1                                                                                     ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��    ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ���$UI_PANEDATA 1(������  	�}/frh/cgtp/doubdev1.stm 8981&action=100                                                                                        )prim                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ��     �N    }/karel/peeritp 1.stm m                                                                                                        )dual                                      }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           ������������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}                                                                                                                               )                                           }                                                                                                                               )                                           )                                           )                                           )                                           )                                           )                                           )                                           )                                           � �����������}�                                                                                                                              )�                                          }�                                                                                                                              )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          )�                                          ��������������$UI_POSTYPE  ������� 	                                    �$UI_QUICKMEN  �������                                  �$UI_RESTORE 1)������  ��                                             �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �$UI_SCREEN ?�������  u1sc  u2sc  u3sc  u4sc  u5sc  u6sc  u7sc  u8sc  �$UI_USERSCRN ?�������  u1ks  u2ks  u3ks  u4ks  u5ks  u6ks  u7ks  u8ks  �$UNDO_CFG *�������      �$UPDATE �������KS_24 �$USER_INFO 1+�������  0%FOLGE011                                    %                                               %                                               %                                               %                                               %                                               %                                               %                                               �$USER_OFFSET .�������                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                          ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                                   
                                        �$USEUFRAME         �   �$USRTOL_ABRT         �    �$USRTOL_ENB         �   �$USRTOL_GRP 1/�������  Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz      Cz  A�  A�  Cz     Cz  A�  A�  Cz     Cz  A�  A�  Cz     �$USRTOL_MENU            �    �$USRTOL_MSK         �    �$USRTOL_NAME %�������%�                                      �$VCCM_CFG 0�������    �$VCMR_GRP 26������               	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                                 	      %~XC56 ****************************            ����            �5   A@  Ap  C�                                                                                                                            	                                           A�  A�  A�      	                                       B���B���    B���             	                                                                	                                      	                                      	                                      	                                                                	                                      	                                     B���                                                    �$VISIONTMOUT        ��  ��$VISION_CFG 7�d��f FR:\VISION\DATA\                   �� MC:\VISION\LOG\                    UD1:\VISION\EXLOG\                  ' B@ �� ��     �                                                                                  �  =	 1- n6  -��         B@         ,             =���=���            MC:\VISION\TRAIN\                       �$VISION_GRP 28������  ( 	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���             	 =���=���=���=���=���=���            �$VLEXE_CFG 9������    1-e            �$VMPHASE  ������          �$VSHIFTMENU 1:������ 
 <�              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ����              %�                                      ���	LIVE/SNAP     %vsflive                               ���VISION SETUP  %vsfmenu                               ����              %�                                      ����$VSHIFT_CFG ;�������	�          %�                                        �5   @   �  @����       A�  B8  B  B�  Ap  Ap  B  A�  B�  B    �  ���������$VSHIFT_MEP        ���   �$VSMO_CFG <������    �z  �$WAITDINEND        �   �    �$WAITDINOK            �    �$WAITDINOUT        �   �    �$WAITDINST        �   �    �$WAITDINTIM       ��   �    �$WAITGINEND        �   �    �$WAITGINOK            �    �$WAITGINOUT        �   �    �$WAITGINST        �   �    �$WAITGINTIM       ��   �    �$WAITRELEASE         �    �$WAITTMOUT        ��  ��$WAIT_ACTIVE         �   �$WAIT_DATA =�������%$FOLGE011........................0006     �$WAIT_RDISP         �    �$WV_AXSRST 2>�������                                  �$WV_GRP_IR  ������ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �$ZABC_GRP 1?������  , 
        2                                 
        2                                 
        2                                 
        2                                �$ZMPCF_G 1@�������  0     
                                              
                                              
                                              
                                         �$ZMP_GRP 1A������  �      � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��        � 	                                     8�                                                     	                                     8�?�              ?�              ?�                   	                                     8�?�              ?�              ?�                   	                                               ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��    ��  ��  ��  ��  ��  ��  �$ZPCFG B�������        �$ZP_CYLINDER 2C�������  �          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                              ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZP_GRP 2D�������  � 
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�   
                                                     	                                      	                                          
                                            �   �A�  �$ZP_SPHERE 2E�������  �      ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                          ,(  ***********************************      (  ***********************************      (  ***********************************                                                                    �$ZZZ         ��    