��   t��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���U�I_CONFIG�_T  d �9$NUM_MENUS  9�* NECTCRE�COVER>CCOLOR_CRR�:EXTSTAT���$TOP>_�IDXCMEM_�LIMIR$D�BGLVL�PO�PUP_MASK��zA  $DUMMY54��ODE�
5CFO�CA �6CPS�)C��g HA�N� � TIME�OU�PIPES�IZE � MW�IN�PANEM;AP�  � � �FAVB ?� 
w$HL�_DIQ�?� qELEM�Z�UR� l� S|s�$HMI��RO+\W AD�ONLY� �T�OUCH�PRO�OMMO#?$��ALAR< �F�ILVEW�	E�NB=%%fC �1"USER:)FC[TN:)WI�� I* _ED�l"V!�_TITL� ~1"COORDF<#/LOCK6%�$F%|�!b"EBFOR�? �"e&
�"�%�!�BA�!j ?�"B�G�%$PM�X�_PKT�"IHE�LP� MER�B�LNK$=ENAB��!? SIPMAN�UA�-4"="�B�EEY?$�=&q!E�Dy#�&UST�OM0 t �$} RT_SPI�D��4C�4*PA�G� ?^DEV�ICE�9SCREVuEF���7N��@$FLAG�@�d&�1  h� 	$PWD_A�CCES� E �8��TC�!�%)$�LABE� 	$	Tz j4@q!�D��	 &USRV�I 1  < �`� �B��APRI�m� U1�@�TRIP�"m�$�$CLA?@ �����A��R��R��$'2 ~����R�	 �,��?���/Q=Q8R3T.Q-R��)P�  1T�w_��
 ��(/�SOFTP�0/G�ENLINK?c�urrent=m�enupage,935,1�_�_�_�_o��Ao/oAoSo eowo�oo�o�o�o�o �o�o+=Oas ������� ��9�K�]�o����� "���ɏۏ������ 5�G�Y�k�}�����0� şן�������C��U�g�y������� TPTX�����:�ٯ�� s �Ƿ���$/so�ftpart/g�enlink?h�elp=/md/;tp�Q.dg��F��X�j�|�5�&�#�pwd2�ɿۿ���4� #�5�G�Y�k�}�ϡ� ���������ϊϜ�1�@C�U�g�yߋ�aT��A�oP��QR�� ($ ����������(����A2QN�PSr_$PS���^�
q�2QR����RU��ʡZ��	���������L�L�Y�S�2 �1�E=PR �\ }mPwREG VED���6�H�wholemod.htm\��singlm�d�oub��tr�ip��brows����I����� ��3EWi{�3��W�i�dev.s�r�l���	1�	t ��	��o� �]�����(/� �@@/R/d/v/��/�/�/�/�/�/�& @</?#?�/G?Y?k? :6+�#//�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O� �O�O#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogo5/�o�o �o�o�o�o 2D ??hzI[��y? �?qo
���)�R�M� _�q����������ݏ ��*�%�7�_W�Q� �������ǟٟ��� �!�3�E�W�i�{��� ����ï�o���"�4� F�X�j�|������Ŀ ֿ��������ͯ f�a�sυϮϩϻ��� ������>�9�K�]� �߁ߓ�a��߭����� ���#�5�G�Y�k�}� ������������� ��Z�l�~������� ���������� 2 hz1�C�)��� ��
)RM _q������ ���/	/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?I� �?�?�?�?�?O"O4O FOXOS|O�O]OoO�O��O�J�$UI_T�OPMENU 1��@QR� 
XQ�1)�*defaul�t�?�=	*le�vel0 *HP #8_& o__m_�Rtpio[23�](tpst[1�X�_�_�_BVX_�_�!$
h58e01�.gifo(	m�enu5Bi9`da1!3BjcbAjad4ikPoa���o�o�o  $6�2�o_q�����Htprim�=dapage,1422,1��� �/�A�Le�w�����譏��N��vclass,5ȏ���!�h3�E�P�܌13L�@��������ʟQ��|53���*�<�N�
Q��|8�������� ��ѯP�����+�=�O��9PQ_��B]�y�aw��oÿ�Vtyx�]�_�Qmf[0�_���	�c[164�W>�59�Xa�oٿ{�]h2�ogm��}j�o sgAk���cg�y�F�X� j�|ߎ�寲������� ����0�B�T�f�x����ۍ2�������� �����O�a�s��� ��&�8�p������� ۟�14�^p���%��sainedi���|%�wintp�p 0bt����6Q r���fo��// 0/B/T/f/x/�/ o�/ �/�/�/�/??,?>? c?�o�?�?�?�?�?�?  �OO)O;OMO_O�? �O�O�O�O�O�O�O~O _%_7_I_[_m_�O�_ �_�_�_�_�_z_o!o 3oEoWoio{o
o�o�o �o�o�o�o�o/A Sew��������o�0���@���⯿]?o��s���������u��d�f� ��&�4����B�h�����6��u7���0� ���'�9��]�o� ��������F�ۯ�����#�5�G�64�1 C���������ɿԯ� ���#�5�G�ֿk�}� �ϡϳ�����2����@�1�C�U�����6\߀�ߣߵ�����4Ӝ74��'�9�K�]�� �����/z������� ���"�G�F���R�|� ��������������p? 1CUgy�Vϯ ����	�? Qcu��(�� ��//�;/M/_/ q/�/�/�/6/�/�/�/ ??%?�/I?[?m?? �?�?2?�?�?�?�?O !O3O�?WOiO{O�O�O �Ol�~��O��l�
_ ._@_R_w_v_�_�__ �_�_�_ooo*o<o No�o�o�o�o�o�o �oHO'9K]o �o������| �#�5�G�Y�k�}�� ����ŏ׏������ 1�C�U�g�y������ ��ӟ���	���-�?� Q�c�u��������ϯ ����O�O;��O�_ ^op���������ʿܿ �\���7�6�H�Z�l� ~ϐϢ�po������� !�3�Eߜ�i�{ߍߟ� ����R�������/� A�S���w����� ��`�����+�=�O� ��s������������� n�'9K]�� ������j� #5GYk&�� ��ϲ�����/ /0/B/�b/`/�/�/ �/�/�/�/�/?��?? Q?c?u?�?�?��?�? �?�?OO�?;OMO_O qO�O�O�O6O�O�O�O __%_�OI_[_m__ �_�_2_�_�_�_�_o !o3o�_Woio{o�o�o �o@o�o�o�o/ �oSew���� z���??*�<� N�`�r���������� ޏ����&�K�J�\� *?������ɟ۟�D �#�5�G�Y�k�}�� ����ůׯ������ 1�C�U�g�y������ ��ӿ���	Ϙ�-�?� Q�c�uχ�ϫϽ��� ����ߔ�)�;�M�_� q߃ߕ�$߹�����������w�t*de�fault�w�*level8ˏ�i�{��7� t?pst[1]�����y��tpio[#23�����u��n����6�H�	menu_7.gifI�
h�13m�z�5��g��e�4��u6m����� %7I��m ����V���!3EW�pr�im=h�page,74,1\��з���pcl?ass,13�/@(/:/L/^/��5d/@�/�/�/�/�/�� �/?.?@?R?d?gy18��?�?�?�?�?�/�6�?%O7OIO[O�mOL��$UI_U�SERVIEW �1�q�qR 
��tON�O�OF�m�O__ %_7_I_�Om__�_�_ �_X_�_�_�_o!o�O .o@oRo�_�o�o�o�o �oxo�o/AS �ow����jo� ��b+�=�O�a�s� �������͏ߏ�����'�9�K��*z�oom^�ZOOM]����ԟ��� 
���.�@�R�d�v���������Я���*maxres��MAXRES�� ����\�n�������G� ȿڿ���ϳ�4�F� X�j�|�'��ϛϭ�� ������0�B���f� xߊߜ߮�Q������� ����'�=�K�߆� ������q����� (�:�L���p������� ��c�������[�$6 HZl���� �{� 2D�� Ucu����� �
/�./@/R/d/v/ /�/�/�/�/�/��/ ??�/N?`?r?�?�? 9?�?�?�?�?OO�? 8OJO\OnO�O#A