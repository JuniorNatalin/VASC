��   �*�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���P�NIO_AN_T�   L $�A* DR  �7SHIFT>V�ALID>I:I�E	IR�&CFG�.� �$V�ERSION �$COMME�NJ �USTOM� @ �2�DE_V_ENB> � �N�TMP�ST�ART_MODE~�NUM_LSJ��� �CHG_�DIG_PR�P�S_MAX���$� ;OP?] MKW>We�STr� ?I_OFS6O�] ��@q�����D<� KDV- KHO�L!�DH*ACT?_INDEX�c!�OPC�o!Kf*Kt)INIT�o �NNOT_NAM�� �$ORDE�= � �#HWl#�"R�EV�(SW1�*2r�*3#� SLO$�� VV3D 8IN��CP16XX_W&C51�D4��C53Y9PKX:PK~�SEARCH�� CHK�TP_�WA� c G�;M�AIN� Q>�2P�ARAM�7EXEyC6�R1SH2�S �HENABL�EpO^#SG_U}O�WD_TI� �;@ C� � P_DoEBUGPBSC,�?CS!DEFAUL�TPB�5�CAPD}U�PWRCLH<�1�KN_IO�A�K��!C�H�F�CFLA�G^#U!P�PWOFF_ALA� �BR� c"DBW@V��0�C.W�C�"2SY�;T[IO� �BOARD_S�!9B�T6�OP�YABD �XP�XMIS�U��W�ALM�Z�W��@`�U>A�Z� �YSM�VH�R� �XDc!iT�[�WmNOP fREAD�0�TS�T�D�fQ�1�j2�j3�UUP�DAT��0RC_�FIN@��aSI�Z�gJD�e>B�eDE��uPTH�fGR�OU��cOUJULONG�!Nt�!NtT1Nt4Kw5Kw6Kw�7Kw8KsBYTE �C�r�C�r1�tvq�t �q�t�q�t�q�t�q�tM9�w10��x1�x�1�x ��x1�x1��x1�x1�2�(��2. (d�f F)@�DI)0�ELTA#���	O�PT��W܆IOR_TRAN��ڄ�!RST�0��a��RESE�^PLI��1�S�"�INT#VL`L&X��O�!d�HO!$@ڀ�`@�ڀ�`@�U@RT�#���#��3�� vq���q���q���q�� �q���������(� ���@��ҙX���8p���FW_���1� 5 ��Wa�cN�CFIR�P@� � &DB. �{ �
BASE�V) � UsI��� vs��vs�료s���s�/�뢈���Y�T��6��~�y�Pb{���o � �RE�@p��>A!5LAYw���bt��}ADD �@�W��W�t3W� �T�5\�6\�7\�8���IA� �� ���!$CNaT��uP�6��RI����PROC�`���` ���`�źB�D ����0�#�5Ϙ|��ǘ� A� �"X0���վ ��TYP������IP: < �����MAS�0��;pT�� ���QMSC�=�� �PrP>�Q�")�چ� O��"�D�!tF�UNK� �F��EXIl�C*`BUSY~���6*`�5��P� �槃@ B� U�Pr�F��FWV��SN��H���X1�`��� ��OCEX� A���� MAC��ML{FB��F_IP-����F_GW3�R3_1&U�U��SàCOU� �Ap�P1�� �� >AX3>A�>At3>Ay� >A��>A��>A��>A���� O�B��O���Z� ��e���p���{����s���s�USX3Oj� Pt3O��O��O��PO��O����L��� � $PA�TH_XDЀA ����	c�� 	c� (u#���N��E�� ����$DOWN�LOA�9@�ARAp܀�#M�" Я���l u����ً������S�NU�K_��&�K8! B�OPER@�8�A��CHE��J!��D$	bhS%�#	cB:�	2A'CPYA%��#LO� ^&�11A'�1�O(SE�R&��A'P ���'��B!��&�&t1�(��eB�K$�@0BUP� Y�5R e&.6�2�'�#7�!7 �"���)���)���)����#�a_BT'#�2DTV�5���3�d�5�6 B!���C�5�C�5�s�5 �s�"�8��D��D�� ,D��@�'�RvG5P���BADb@�WNGsGS�G$�TIN:`N�EAFE��@_��&��LD�9I�A=���P���P��SERVLI,�(�h!o���{���#CM:WSVFZLOIW	b��fW��NR���'IO5��V곐�в�pU�U��"�~dMOn�b$H!CM� �S��b�@t�NY�e a#c�tet�.f+�D&d�CLzf0�_+���ID _� [�lge�lg o�lg��lg��lg��ްYNC_�vc�e�c �bsf�e�k�c�e�c�e��c�e�cHp� L�1v��C!C! �s!�s!�s!�s! �s!�s!�Nr�Nr|Rw(�CLASS�`[����ve���؏��L� 	 � }ΪENABL����ES��+PENG�THJ>��_�UB09������DA7�S��]�ϠR�ERRDE�AC�I#�NDEX��3p���VPaQ�b�h��IM0x
�� $��H�"��L"��ET���V�񇠉Hٰ�bR5�0�B�F�"I#�����R_�N`P QIALB�$R7�0<Q1���$VMA��M.TSIMS��El���" ���AƠ � 
Ϊ9���>�㤽��PU%�摝��� ��]�_�4���WRKxH 1v;v��	���`�0�"�\�TP_DEBUG�"гO�_�GPWO*0"�!W�  �a�Ns�������ɥ��OM����UBcYT�����$S_�SYSY����U�g�y��ϝ��$�s  ������Y�a �N��#AN 2 ���N� &�� ���������Խ�ǲ��ǲ$�ǲ
-�ǲE�ǲA]�ǲȰwϽ���ǲ��ǲ��ǲ��$�Ͻ���ǲ�ǲI�ǲ 5�ǲ"Mߒǲ$e�w�&}�w�($��w�*��w�,��w҉.��w�0�߂��"C�FG ���V820P02 ?131028����a��O���P���� ���� �~�wЀś�@�����X�� X�F�ANUC Rob�ot Contr�ollerC�A�05B-2600O-J93 ��V|��� �  X!�Y� ��Y�dm�=������G ����U���, ⿱e���f�m�c:pniotrc.txtX�����X������=�2 "�L�@B�&��N�C�y���Sװ����). �b��� 2�� h�CP1604 �DAP V2.6Hi�L�!"�X�#"��p�%"���'"���5�"��7"�)"� �1�m�L�� "�(M�����������16����+=Oay�����
�XX{i���/"/� O/�/�/�/�/?%? 7?I?[???�?�?�?��?���������?O(O�?I���G ��!� .1.���tM�1� ۝<۟<tO7OID����� �kj�ltvl4116�30r01rs--kux�O	__-_?_Q_���V_z_�_�_�_�_�__WS7-PC�_oo,o>oPo boe_�o�o�o�o�o�o��j!172.26.29.17hO�c255.&u�bx6��=Z~� c�������� &��m6�Z�C�~�m� ����Ə���ُ�VN u�) � �!�Y�k�}��������ş�=L ��A�MC:PCST_1.X� ��+��AUD1:\P�N2610.FW_L 3.9J�l+��i����Xd )d����������� ʯܯ� ��jo6�H��Z�l�~�����7�FR:S7PRJ��ֿ�9���\fw�_image.fwW�!�.�U�g�y�>�� ,X����h�|��@n ���H��@��C����� x���e�e�g���EE?E�����(�*�z (g��^!!����7�d�r	y�>��ST 2	�J��YD{?5�?������ p?����"������E�J��!��K�5�@��Y��*���콟��!�m��������"� �U���H��1�i��G�Y�k������  AJn��������sA�2�e�҄�
> y�K�o����ۅ�xԱB�1��b ���#5G�w
���xԲ���������/+��\3/E/ ?�xԬ�t/�/��ܞ(U�/�/ ���ѥ!e/�/? �&8C?�?�? F߼?�?�?�?O(O:O 	O^OpO�OQO�O�O�O �O�O _�O$_6_H__ l_~_�___�_�_�_�_ �_o�_ oDoVo%ozo �o�omo�o�o�o�o
 .�oRd3�� �{�����*� <��`�r�A������� ��ޏ���я&�8�J� �n�����a���ȟ�� ����ߟ4�F�X�'� |�����o�į֯��� ���B�T�f�5��� ����}�ҿ���ſ� ,���P�b�t�CϘϪ� �ϋ��������(�:� 	�L�p߂�Qߦ߸��� ���� ����6�H�Z� )�~��_������� ��� ���D�V�h�7� ����m���������
 .��RdvE� ������* <`r�S�� ���/�/8/J/ /n/�/�/a/�/�/�/ �/�/?"?�/F?X?'? |?�?�?o?�?�?�?�? OO0O�?TOfO5OxO �O�O}O�O�O�O�O_ ,_>__b_t_�_U_�_ �_�_�_�_o�_(o:o Loopo�o�oco�o�o �o�o �o6HZ )~��q��� �� ��D�V�h�7� �������ԏ���Ǐ �.���@�d�v�E��� ����������՟*� <�N��r���S����� ̯������8�J� \�+�����a���ȿڿ �����"��F�X�j� 9ώϠϲρ����Ϸ� ��0���T�f�x�G� �߮��ߏ�������� ,�>��b�t��U�� �����������:� L��p�����c����� ���� $��HZ )l��q��� � 2Vhz I������ /./@//d/v/�/W/ �/�/�/�/�/?�/*? <?N??r?�?�?e?�? �?�?�?OO�?8OJO \O+O�O�O�OsO�O�O �O�O_"_�O4_X_j_ 9_�_�_�_�_�_�_�_ �_o0oBoofoxoGo �o�o�o�o�o�o�o ,>Pt�U� �������:� L�^�-�������u�ʏ ܏�� ��$��H�Z� l�;���������؟� ���� �2��V�h�z� I�����¯�����
� ٯ.�@��d�v���W� ����п������� <�N��`τϖ�eϺ� ���ϭ���&���J� \�n�=ߒߤ�s����� �߻��"�4��X�j� |�K���������� ���0�B��f�x��� Y������������� ,>Pt��g �����( L^-���u� ���/$/6//Z/ l/;/�/�/�/�/�/�/ �/�/ ?2?D??h?z? I?�?�?�?�?�?�?
O �?.O@ORO!OvO�O�O iO�O�O�O�O__�O <_N_`_/_�_�_�_w_ �_�_�_�_o&o�_Jo \ono=o�o�o�o�o�o �o�o�o"4Xj |K������ ��0�B��T�x��� Y�����ҏ������ �>�P�b�1�����g� ��Ο������(��� L�^�p�?�����u��� ܯ��$�6��Z� l�~�M�����ƿ��� ��˿ �2�D��h�z� ��[ϰ����ϣ���
� ���@�R�!�v߈ߚ� i߾����߱���*� ��N�`�/����w� ��������&�8�� \�n�=����������� ������"4Fj |�]����� �0BT#x���k�$PNIO�_IM0 
�����N��k� V�A05�B-2600-J�930eF1�73� ��k���LST 2�	�Dn;*�?�e�F'_$g|/K#�`R(�b/�/B+�$bY!�/�/�/��(��/�/
??�54�PZ/8?�?L"�y4�j?|?�?�"��$�1�#�!��?O�?�1�/OO �$�1)3�?�OC+��D��?�O�O"H 6D�A�?�O�O�K9O_)_  J�H)?[_m_ ?�T��O�_�_
"X�P
�T�/�_�_Po	_7oA-�ed��_(ho�o"b�`�do@�o�o�o]oA-�1t!��o4��"FTeq %{��{I_��&� ]8�\�n�=������� ��ڏ���͏"�4�F� �j�|�K�����ğ�� ����۟0�B�T�#� x���Y�����ү���� ���>�P�b�1��� ����y�ο࿯��� (���L�^�p�?ϔϦ� �χ����Ͻ� �$�6� �Z�l�~�Mߢߴ��� ���������2�D�� h�z��[������� ��
����@�R�!�d� ����i��������� *��N`rA� �w����& 8\n�O�� �����"/4/F/ /j/|/�/]/�/�/�/ �/�/?�/0?B?T?#? x?�?�?k?�?�?�?�? OO�?,OPObO1O�O �O�OyO�O�O�O�O_ (_:_	_^_p_?_�_�_ �_�_�_�_ o�_$o6o Hoolo~oMo�o�o�o �o�o�o�o2DV %z��m��� �
���@�R�d�3� ������{�Џ⏱�� �*���N�`�r�A��� ������ޟ��џ&� 8��\�n���O����� ȯ������߯4�F� �X�|���]���Ŀֿ �������B�T�f� 5ϊϜ�k������ϳ� ��,���P�b�t�C� �ߪ�y߼�������� (�:�	�^�p��Q�� ������� ���$�6� H��l�~���_����� �������� DV %z��m��� �
.�Rd3 ���{���� /*/<//`/r/A/�/ �/�/�/�/�/?�/&? 8?J??n?�?�?a?�? �?�?�?�?O�?4OFO XO'O|O�O�OoO�O�O �O�O__�OB_T_f_ 5_�_�_�_}_�_�_�_ �_o,o�_PobotoCo �o�o�o�o�o�o�o (:	Lp�Q� ���� ���6� H�Z�)�~���_���Ə ؏����� ��D�V� h�7�����m���ԟ� ��
��.���R�d�v� E������������ï �*�<��`�r���S� ����̿����ѿ� 8�J��nπϒ�a϶� ���ϩ����"���F� X�'�|ߎߠ�o����� �߷���0���T�f� 5�x���}������� ���,�>��b�t��� U������������� (:Lp��c ���� �6 HZ)~��q� ���/ /�D/V/ h/7/�/�/�//�/�/ �/�/?.?�/@?d?v? E?�?�?�?�?�?�?O �?*O<ONOOrO�OSO �O�O�O�O�O__�O 8_J_\_+_�_�_a_�_ �_�_�_�_o"o�_Fo Xojo9o�o�o�o�o�o �o�o0�oTf xG������ ��,�>��b�t��� U�����Ώ����� �:�L��p�����c� ��ʟܟ�� ��$�� H�Z�)�l�����q�Ư د꯹�� �2��V� h�z�I������Կ� ��ǿ�.�@��d�v� ��WϬϾύ������ ��*�<�N��r߄ߖ� eߺ����߭����� 8�J�\�+����s� ��������"���4� X�j�9����������� ������0Bf xG������ �,>Pt� U�����// �:/L/^/-/�/�/�/ u/�/�/�/ ??$?�/ H?Z?l?;?�?�?�?�? �?�?�?�? O2OOVO hOzOIO�O�O�O�O�O �O
_�O._@__d_v_ �_W_�_�_�_�_�_o�o�P�$PNIO�_MOD 2����;aN��  @DAP V2.6o��Phdj`ka�_�SAFE 8 B�YTEzohc�hd{o32�o�V"hd7hc�fka �o~hdUa�d�b�as ^p�_����� ���$�6�	�Z�l� ?���������؏ꏽ� � �2��V�h�;�z� ������ԟ���˟��.��R�d�v�+gST�M  ;eNja+q����Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T��f�x���O_WR�K ;i ���_j�bC��� p��	�