��  	��A��*SYST�EM*��V8.2�306 4/2�
 014 A�5  ����A�AVM_WRK_�T  � �$EXPOSUR�E  $CAMCLBDAT@ �$PS_TR�GVT��$X� aHZgDIUSfWgPgRg�LENS_CEN�T_X�YgyO�Rf   $C�MP_GC_�U�TNUMAPRE_MAST_C�� 	�GRV_}M{$NEW���	STAT_R�UNARES_E=R�VTCP6� %aTC32:dXSM�&&�#�END!ORGBK!SM��3!�UPD��ABS�; � P/   $PARA� �  D��ALRM_REC�OV�  � A�LM"ENB���&ON&! MDG�/ 0 $DEBUG1AI"d�R$3AO� TYPsE �9!_IF�� D $ENwABL@$L�T P d�#U�%Kx!;MA�$LI"��
i�8�APC�OUPLED�� $!PP_PR�OCES0s!�(1Ns!���!> Q�� � $SO{FT�T_ID�"�TOTAL_EQfs $0'0NO*2�U SPI_IND�E]?5X�"SCREEN_NAMr {�"SIGNe0��/�+!0PK_F�I� 	$TH{KY�7PANE24� � DUMMYE1d�4d!�54�1�@�ARG�R�� � $T{IT�!$I�� N DdDd D�0DU5�66�67�68�69�70�7G�1EG��1E0G1:G1DG1�NG1XG2cB��ASBN_CF>"� 8F CNV_�J� ; �"L A_C�MNT�$FL�AGS]�CHE�C�8 � ELLS�ETUP 	 �P� HOME_I�Oz0� %5SMA�CROARREPRJX{0D+>0�dR{�lT��AUTOB�ACKU�
� �)DEVIC&�3TIc0�� 0�#��PBS$IN�TERVALO#I?SP_UNI��P�_DO�V7�YFR3_F\0AINz1���1�S�C_WAx�T�Q-jOFF_� �N�DELZhLO�G�R�1ea�R?�Qf`�3?�� {1�5��h�MO� ZcE' D [MZc����aREV�BI�L�g�AXI�� �bR  �� OD7P�a�$NO�@M�#��cr�"w0� u<q��`Z0�D�C d ^E RD_E�`Ts �$FSSBn&$�CHKBD_SE��UAG G�0 $SLOT_��V2�q� Vzd�%{���Q_EDIm   � cQ�G�CPS:`a4%�$EP1T1$O�P^02dap_O�KnrUS�!P_C�� �q�T�vU UPLACI4!TQ?��p( ��QCOMM� e0$D;�Q�J0f`�y�?��24�BL%0OU�r ,K�QQ2$QU B�@y O]Åޗ�CFWt ?X $GR� ���MBZ`NFLIx���0UIRE���$g"� SWITC�H��AX_N)PS�s"CF_�G�� � 
$WAR�NM"`#!�!�p�@L�I�f�NST� C�OR-�RFLT�R`�TRAT;PT|b�� $ACC�Q�N ��r$OR�I�o"�RTlP_�SFg
 �CHUGz0I��bT��1�IʐT�	���K�� x� i#
Qnr�HDER�2J; �3I�2D�Q3D� F�5D�6D��7D�8D�9s! ���CO�D <�F �����#�܀O�_M�� t� 	PEq0�1NG�1iBA� Q���q ��!�Qp�0=q�0�I�P�PJ�t�G�S��pm �RC ��4���"J��_R��g�C��J����ļJVep�%C�X���p0�h l�AzOF�� 0  @F RO0��&9�6�IT3c9��NOM_yV�lS� $��D Ԁ0��A�B�'&�EX��B0��P����
$TF�E0��DM3N�TO�S3U8P�+� -0P_H��j 1�E{� �%�Y#&�d%(��1��$�DBGDE}!m_p$��PU��1a2)��I"���AX�Ae$]eTAI.�SBUFivX�/� � k�f�P�I�$��P��M���M��^���F��S�IMQ� �$K;EE:�PAT0������N#��Y"�$�L6/4FIX/���&�TC_��� ���c��CI됎�PCHOP��ADD���� �����I"m0p�3�_��!f���n!
��a���W���d"@$�M�C�� �0yJB�E�ͤz��l�+�i� sTN��� ��p�CH� EMP�#$G�����p_�lS��1_FPm��@��SPE��lPn�������� V�q<r�A̛�JR�<rSE�GFRA��3 �R>�0T_LIN{sMPVFs!�$�'�_�"�#m�"� R��D$�y� D ) ���`�����2�f��)P���Ţq�f�SCIZc��T����3�RSINF��G�R �e3 e��> L�з�ΚCRC(�AcCC n��3 ���*���1Ma�������D&�e#
)C+e`T�AM ^�&�T(E�VT&i�Fj!_F��N�&�@f�`�((�������'� rj1���A! �>p���-�RGB�ª�F�B ׂ��De�R��LEWر�Q���<�/�. ���Xs"� ��Ư��5b�#�R� HANC�$LG~��!�Q U�y�gp��6�A:`� a�c�R?2 �3p0���3\��8RAnS�3A�Z��7HP ��O�F#CTC�Y07�F)�����R�ADI�KO �H@�@�o��D~�.��6�S�p����qCMPW*���M�4GAES��l#���0�I_�4#  z�I+$�CSX���H���$*�?p�s��T��B�C�0N�p�I�MG_HEIGH�mqrSWIDK��V�T��M��pF_Ap {��B`EXP�A�4��U�CU7�]�U�%�% $_�TIT&���r�s�p��LE:RZ_% {�&*��{� ��A~�NOwPAD	q?W�i?�,����x�DBPX�WO�&�'��$S�K���r Y�`T�0TRL%�( ��,�A!���@��rD�J��LAY_CA�L�q	��`�@�gPL�	�G�SERVED W�wb�w��'��T	���9��0����`dAA%�)�b��PR�? 
��D"����%�* _���$��$"��L2oy+|"Ѹ��&�y,�"��PC%��-�"�8�PEN�E���!.�"�4�OqRE}��r/H��0C�� *$L2�+$os��+@C�hT ��O�0_D�A��RO�����|��|�RIGGE𞖄PAUS��VE�TURN���MR-_�TU>��a��EWMF��GNA9L����$LA-���n�,$P��-3$P\@!�.�b�b�C!�!��DO` ���\�H��b�GO_oAWAY8�MOD��0�B��DCS�rpEVIm� 0� P $іRB��
�PI���SP=O��I_BYT2��ҽ�TXw�L$�1 �H� 7��Ф�TOFB��FEl����إ�w�CU2�DO����0MC��N���P7�`����Hy@W�� �w�ELE�GR3 T����cCI�NKh�����U�LƘ�HA����$<���� ,w���4 ��`MDL��� 23��(�O��^����C�2����J]�}O�m�}2�@U�r�h�������	��溥@w�%U5� $]��0�PcC�P@Z��Pa5бw��ϲ��̵IDJ�˶�b˶9W ���NTV��в�VE��(РW�D�2�W��J�&���pS�AFE)���_SV>�BEXCLU�a���>2ONL���Y�6��3x@�Qw�I_V|�@�PPLY_����� Ƕ��_M�">��VRFY_�c��	MS3�PO��x@!֧@1~S4�^�O���İ���@� 6��`T�A_ ����  � ���SG�  w7 ��CURπ��}S��tpUQO�REaV�ٯҦ�jPUN�p@��ԥ��Ё������0���ѧ@���  Ӹ��PаI�r8 �@� F���T�OT �At<�At'qAt^�� `+�M��NI>�r9 L �`���Aʱ��DAY	�LOAD��6tv�zBs5>q�EF�P�$�X�:�' SO�������`_RT�RQX�; D�!O��RQ{������:| C7 �D��A;`���< 0��Z��p�Z�>��6DiU5��bCA��g =9�[`NSk�6��ID� PW93U�4���V��V_U���< �DIAG�r�u>8 *$	V��T%ep�
p�R�r��{Vn2`��SWB@��u���R ��;��f �OH�r�PP2a&�IR�Q�B����m�����|	�BA ����D@�������=��CY �RQ�DW�MS� A�Z`w0{LIFE �`�/Hq��NB��K��@��!����CV�@f�NЀY0΍QFLA�4��OV�@W.`�NSUP�PO�`�A���`_���z_X�C�a�
�Z�W��A��B�8��CT%U? }`��CACHE�'�C"ۣ�կ���� SU7FFI�ϰ�`�%a6t��Bs6>q �D�DMSW%U@� 8��KEYIMAG��TMF�C�!�с�&INPU}R wh�G�VIEL �1A �BGL�/đ��?� 	 �`PfPcBMP�!g�1IN^�Tb��	UBFv�JB�a�d��O#Q	T�3��S��Uu59d^�;8�OF��H���C �Va!gOT�F��ץ1�D[�P_GAI�Q���@�@̒��NI_�0C���5����6�PTIC��O �PE���"��}1�A{��PCF�@INy��P[E�Aq�@!����A$P�3D  TP��6D�7I�8T�r=�Rv�=�AVE�F�FBP�c�C���3AW_�@<���E���v�DO<4SLO��>�1TERCE/���bDL/`�J3UFU' RQ�E�e{0�P�E}1�D/��B�FE��3 N��3qPQ;`�5�R�6��R�5@�G�FF� 䠣�$�p1��G �1�0���1F ����0�3�0 ��AbyB��cCARRg#i0�9T$ <2%cyftqcRD_4�06FSN�����T� �FSY��D�I"e�C��A�DĔ�dEG�R�F #	X2u0��Hb�C9 �0ǰY���1�@3��G  �2A I� { _��3]6�0�s�1�s�1�r ���D Ц$J�z�STp@!�r)��tk���tv��t���pEMAaI���/1� SB�@AUL��K�")8}1�COUdP��P�sDT!���L,�@d�M�SU��ITh��RZ�U'}�N��F SUBRT��C봅��*rw�SAV~�@� �ES��m�������P���M�ORDM�p_pRPd���ډOTT���A��P�60��s��#AX��,��XRP���DYN_�B>�Mb��6� ����G3��@IF� ����b=�N�� �05��r�C_RO�IK�"���҄���@R�!���8��D�SP�&��PA��I (v���ß���U���5D��M�pIP0Á��D  ڔTHR#ES�`˕��TZۓHS�bۓR`�E[@��V����@�㑤P��NV��G����]�ؖRPFB��d���@(�F�!SCbRu��M-P>��FBCMP�À��ET�a��O�"FU��DU'��QPPEP���CDљ[���-3��� NOAUT5O��P�$z���z���PSy�CR��C�BE  �8v����QH��в ��r�г���@N��� �S��k���v�������T�!��7��8��9���B���1�1�1�*�17�1D�1Q�1*^�1k�2y�2��U2�2*�27�2D�U2Q�2^�2k�3yʥ3�3��3*�3�7�3D�3Q�3^�3�k�4y� 
 v�O�UT� ��R � �"@	WvPRuPLC�WAR+v�`����R|�$FACm��SE��$PARM1��2m�"k����x³�pA l��EXT��!S <�)9I�g�0Rv�������P�FDR~dTT @  ����E-�BE�11N(OVM�4T�A\�oTROV\�DT��|�MX��vP&�{�N��IND��:
���`E�PG3���� pb1�`DRI�@�cNGEAR�1I%OQ�KL��N�@:EFF\�k�� ���Z_MCM1�E��F�UR5�U y,��V�? �F0@?� Ð0�yEi@� ��p���2� V�RTP��$VARI�5�����UP2_ 3W *�?�TDI�iA�>�TV��  �x�BACG�X �T�p@�U�=0)$/PROGC%?���:�b�IFI�� �wYPa��!@��FMR2�Y ,�k��B-�Mp� 1�8J\s�}0p�L��_���AC@IT_<[U�C_LM��>(DGCLF����DYt(LD���5�������T��uZ,&) � S؀�t�[ P�P�":2��$EX_�!�(�!1P'�נ���!3;56s�G���\ ���2��4l�ON����1��T�1Q�GR��Un��BKU�O1��7 ��PO��9Є0$�W5�0M6`LOYO��1SMw`E��������`_E �] ��V�����,PM�5^�5���ORIp�1_�5O?L �SM_M	r�0`�5R��TA/I�a�5XPO�UP�:P b� -���b]$�5v@^r��G{J� ELT)@��AUS�@ONFIG��A� c1aCrD�_$U+aא$`}��A�@P� OT�G���TAk�-�3SNSTv`PAT`�f`ROPTHJ(�N�E� 8��W��BARTE`�E�p���r�AR[pRY��SHFTR��AQCX_SHOR1�K�.F% 9@$HG�Pa>!.�GOVR����PItP�;$U�� M�AYLO0�!A��`� ��Q8]���]�ERV��Q ���Z���Gv`QR��t�;e��tRC���A�SYMt����AWJ�G����E�?QkibQ�U�d@A�CU�qP��YUP��Pġ�VOR@M�l?0�1 �c�r�2�6P�@!s���q�%d Ƚ��xLTOC�A|�1i$OPo�"����2��pH�O,��Z�REbpRأ��X)�K�ReipRU�u}x[QDe$PW�R	 IM�ubR_�Xs8TVIS/@�b��,r�B e� �$HC!�ADDR�H�1GR/�$���˱R3�����f H��S��N���\��Ӏ\��\�*Â�N�U�o��HS[�MN�!?g uB�trq�[�OL1��h�x��^��0ACRO�p<�AhqND_C1�|�xa�tšROUP���!r_ÐI1�Uq"q1 ��6�2��<���<�Q�=��<�*�<�7�6�AMC��IO��D7�䩓G�t�� �h $� Pp_D��0��ޣ�PRM_+� �,�HTTP_�|�H#�i (=�O�BJE���t$��LES��ְjrN0���AB_���T�3P�S����DB�GLV1�$KRL~�yHITCOU@�Z�1Gf�LOC�O�TEMPt�����zp�v{pSS��I��HQWe��A#�kW��`�INCPU���pIO�e���r������*�IBGN��$l���� WA	I�s�aP����R��ӳFW	 ېLO`m��s|���y�AN�A$Bo��������������RTN/`�CU?F_DATA�㖠����_MG�2/ F��>�S(SE��r��8R�EC���N�b��2�h�I� m )@� N�_h�Y�3tĎH�EXEwɒ�Ф K`_�Xu�0�n�$SCH�`�Q�P�R��FLGvQ #2�	/�oo�����v ��OPÒ�1�~�TRA�B��CS����9�px ;$C�CTA���'�IGN�MoO҈0�M~�Tֈ��v����vN_PCSO8�QUp��ECFBa�� Q���u��Ғ�	\r��aL�������@DFRs8������SPT �$���SEQ_� Z3NS��H�*�ɀ��rC�q�@Xl�SL�}P r�Q �-@o�bc��0��se:!D�IOL]N4q 8��R��$SL�$I�NPUT_�$��p��P- ��d��S�L���!rr��#� yp��ݐF_AS�"s:$LO$�O���Р�r+�����PHqYP���^�  8�sUOR��#t `J� ��(�%�s�%�|���pP�s������|������DAUJR�u �� N��UJO�G�G$DI,�$�J7�dJ8O	7�60I�AXj7_L�ABQHpZ �NA7PHI� QY�=D� J7J8�0�_KEY� k�K)�L�%v  ��AVއP�CTR�eS�FLAG:2��$�LG�$w �����Y3LG_SIZJ��0>� =A�=FDHI<S�1 J;@=:tsC� � �A�j�@��X_R�������5���LNCH2x�����U01#��!BpU��)!(�L2#("DAUN%EA�)�Dtd"�Z GHEr @��M�BOOQ�yt3 Bd��pIT�Ø$p{�e�#ү(SCR���`�D��[2$�MARGI�D�,�X�ctH2��M�S0�L�W�$�M�=$X�JGMC7MgNCH�M�FN�bF6Kl7q�j9UFx8��Px8n�x8HL�9STPx:Vx8àx8� x8RS�9H�`�;U�C�T�3�bX�p7CIU䑌47�R,6� +�22G\9lPPO�G�:0�%�3�d2OCG�{8,���GUIj5I�3�B(3S43Sh0l1��P�rC9��&�P�!N݁-�ANAM�Qq�Q�VAI� �CLEkARfDn�HId��~Sr�~RO�XO�WS	I�W�XS�X8lҸ��i�i1��Tքn�DE�V��,X�!_BU�FFqz� �pT60R$IEM�����'  �
bjqq{�� �p���ˁIpO�S1je2je3ja �P
b~Q	p| �! ߈�aZS��{���IDXtPK�@z�TjK�T��Re Y��~�a {$Ev�C{T��v)v y�ch�} L� s�����������w3���u�Kc�#_ ~ � +�#��!޸s��MC"{ �! CLDP��>vUTRQLI� wT 2 �y�t�����p͑�"nQD��ڠL���t�ORG2 B!��'��������!���s͔� ����tE|�t�SV_PT�p腔R�ǄφRCL�MC݄m��� ���MISC�� d%!�aRQ�����DSTB��` 1K��!X�AXvR� |[�t�EXCESm/ ,-�M���q���?�vT 
 -�T�㠃�M�_��I�����r�����MK�� \�PǻMBۢLICL�B�� QUIRE,CM�O>�ON�DEBU>����ML�������e�H�Pށ�l��2�Di $D�$U�PyACKED����DPxv���IN�b$q�_ Q �pI�U������� ��/�	�=�U�4�T�I���P�MND:!S�Sb�#""$��DC��6$IN]�3'RSMD ���PNr�BCv��y�PST���� 4q�;��fR�Il �e�eANGܭbI�p��AQz���;�$ON,"�MFqT��i���00�uz� 3�SUP~�� ��FX&��IGG�! � �ဃs��#�s6F�tR{�v��b�ɵ��ȵ�x����+�DATA����ETI8 ,�x�1�1`INb� tV?�MD?�In!)M���YӇ�U�H#�SX��DIA!Y�ANSAWe�Y�Pa�AX�Dl#�)@1�ŀ���[ ��CUSV����I�T���LO�f �������G�����5����� � ���MRR22��O� ��J!Á� d$CALI�Q��GrQD�2f`RsIN�0G�<$RR��SW0�����AB�CS�D_J2SE�e�I�L�_J3��
���1SPm I�P�����3���ѓ�I�B��J����āOa�IM��CSKP �z<�- kS<�Jm!��Q<�m�S�m�c��_cAZ˂	��ELa<���OCMP&������1�� ���`1����� ��Z��D�OINTEVpSb����2I��Vp_N²��7�a��43̒�A	DI������DH��6 ���Y`$VQ঳�a$l1$ �!�`��Q$-�2��H �$BE��|�	�qACCEL������ IRC_9R-��ONT�a�c�$PS���rL  �!�s -!sPPATH�	Z�"Z3)����_ga����ʂ�C��� _{MG�Q$DD�<�"$FW5�1�`�����DE��PPABN1ROTSPEE�ka/8�pc�kaDEFۑ�~)$USE_P�J>SP�C�@>SY
 �� ʁ �aYN1�A�c�x&,�o�x!MOUf�NGtB�OLJ�$INC�� ����X��'3�Y�ENCS�P��I�!�V�IN�bI)52��c��VE� H�*223_�U>��<3LOWL��Qz@���p�%\6D�]@I�3� �p�%�C�' #6MOS�P�M�O���`ʇPERC7H  y3OVp t" �7�a�3��_2����� ��b%��P*�A)EL=T*��)�$5��_:�ZFu6TRK�4�bAY��Cܑ�A)�E�C8!��`�RTI���"�`MOM�BX�ܒc���G��D��C\jb� DU2��S_BCKLSH_C) U� �6�0�#��:T�"xEZ�!e�CLAL2`�"2���@�`wUCHKt�p�eS� RTY��B�5$�U�0�_�cN�4_UM���YC�SήSCL�T# LMT��_Lg����T�gE m!`k�Pe���0Q�!&@bd�8P	C�1�8H�pl���U�C뀎rXT� �C�N__�N���f�S	F��9Vb""�7�p�a)u�hCAT�^SHo�_���&U�Q�6��*����PAL�T�"_P�U�C_�p��P�F�0�q�C�t�UJaG�����sJ0OG�g>�BTORQUT �� �3�I�/��2�A��_W�E�D��7���6��6�I>�IL�I�F9�)��#��VC� 0R�J���1ಎ��Əc���JRK������DBL_�SM�!5BM��_D9L�5BGRV=�6�0�6���H_���]d�COSq��@q�LN��������� ��� ��h�Қ�����Z���6�MY���}��TH��1�THET=0e5NK23�[�l���CB`�CB�CT�ASƱ��h������`�SB���k�'GTSE�#!C�� ����|s���ϓ$DU�P>G�D��!����3��AQ��&�$NE�B��I��#���L$~ O�AS�|���c�n�n�LPHq�Z�45Z�S��ͳ��ͳϕZ�ޖP�����~ V��V��T� ��VźVһV�UV�V��V
�V�H�����µ�:q��һUH�H�H��H
�UH�O��O��OI٪��OźOһO�O��O��O
�O��F�Z��������ԑ�SPBALANCE��~aLEȠH_S�S�P��4���4�ϖPFULC8�_�G�_��ϕ!
1���UTOy_�P�uT1T2���2N�Quc���O@�Aa�?�0��ATK@�O���'�INSE9Gu~1REVB�~0�1DIFtEF	1�l+�r1�IPOB!�gQ@��G2����Q�?LCHWAR
"g"�AB�q�E$ME�CH�� ��!��VAX�APEd��u�� �� 
����5ROB�0CR)���b� l�MSK_|��� P ��_R R���+:!vD1r/0-"+ ,3ET+ ��IN��MT�COM_C��� ��  �3� !�$NORE3���OPWO��� �w, k SBU఍�QOP� �T��
U�=PRUN,q�PAR D���\��0_OU�!��S�AB�"$ I�MAGVQ( B�Pf�IM� BIN'��BRGOVRD<��	@P!Ap�!_��q��R�`R�B�`��[aMC_�EDT_� K`N�l�M�JaPMY1�9Ia��nSL�6�" � x $�OVSL��SDI0DEX�c&�cKA "V�!$N'!� 5 %#:'5(��Q3��q_� �" � @!��l"���2� �2
&_����'�!�! `��0�ECT�  �� H(��PATU�SP{@CD�ZD�X�&BTM�'�!I�	�4Ia�#�" � D( E"�"Z�yE4��!FILEJ@gP�!EXE� �Q�72K24t#�{ ) � �UPDATZ1$T�HXNDP�������9T�PG��UB�!���!��!�#JMPWAI2'pP*#�5LO`��F�p�!�RCV?FAIL_C�A��1R�@� �V�a�d��<E�R_PL�#D�BTB�q�UBWDd.F� U�P/EIG8I��TNL#p0D�BRT�� ERV�E�c�D�bD�1D�EFSP�P � L( ���@``�qp�CUNI"7�@�1�RR0!�.�_L�P~�!  d�Pr !� 0�q�!] �ATA$�uNP�K�ET$R#�BUtPsIPB!� h�?ARSIZEp@hE0GQ�RS� OR�#?FORMAT��uDcCO�Q�EM���TSUX� :"p��PLIpB!� � $| P_S3WIp��S0���U@�p@AL_ � �$�AAVB���C�VD	$EZ1��`C_zA� � � Q�Va�J3��V80RTI�A4hi5hi6VMOMENTtc�c�ch�c�c| B @ADtc��f�c�f�cPU��N�R�d�e�c�e�b���S�P H$PIQ��6�H�Z� l�~���!ڦ������� ��GQ�&SPEED�G�R�tE�D�v �DE�,@�v��x�8�y�ESAM#���F��wL�EMOV_AXI�!�z��%����7�z��@1d��2dR	 md��	`a ���INڌ	`/�����؄B�#���#�C�G�AMM��A��R��GET�rFIMS�PDczd
��LIBR�1�BI�@bS$HIB�0_^� f��E`bŘA���ӖLW��  ����$�Ӗ?b���@�aCfEq�|�  $PDCK�D���_.��Pdւ SiaɅ���c���f��~c �$I� R��DW��1"D��LEa�q�!�?h�}�VpMSWFL1D]M`SCR�86��37+�U��qi�q$�S]�p�P��3URB���GR���S_SAVE_DX����3NOC`C�! �2Dd����Sj<v幾 Uy�mp����pW�v(<Ƚ�.aO�AA��� ������e�x��vv���ǜ�ZÌ��1 �rMu� � ��YL5s~�ɇ��~� ����NB�KA���!WѰ�(��4��`������M��L�CLHK�aD�^�1j����PM�� � ό $���$W�Є�NG1]a�� d��#d��*d��1dV@@��s���S��	`XP	O+caZ&��P@tG� p�| ��Uv������,�;�Ca_�� |�Si���i ��c��c��mj	���b�jE@�� ��Jy�� ^`��P�Q��PM4 QUP� /� 88PQ��n�QTH� HO��n��HYS�PES�����UEr�hP��� � 6B;Q#��#��_� 'Ѵt����EN/	PBG _@B�[mB?�#*#�Jہ��I��pEW �vGTF-b"��PO�4�   1�𮗫"UN� Nя �{ �rp� PD�E��-3�B�ROGRA�!�2064M ��ITh@��{ INFO�� �� ������ (v�SL�EQ�v6�u6��${ �D�0p�����QOv����#��E��sNU��AUT���COPY���0��qʰM��N��^��PRU���� gQR�GADJv!�wRX'��B$P&3�&W(P(��$�s	 ��3EXF@YC���!NS�T�; �4ALGOk�.`�NYQ_FREQ���U �w�!�T�LA�hC�!��b.��5CR1E�0��l�IFQq��NAT�%�$_GhCSTAT�@4��M@R���31	���Q�31��|$ELE�0 ��Nb�SEASIr1���"�a2�1�� �6BƀIa�"�q��M���2AB�Q/`E�� �pVU1�6BAS9b�5����U�@� ��g$�1F�|$���� X �2 2� 	����@QFBPGQ|р�eEF|F g~"PFe1=�=GRID��S�B|P�wTYs3�`�| OTO �1Q� �_4!E �BwsRO$��$� ���;LI:�PORAS�C\'v�BSRV0)T6VDI�PT_�p6P�HT��RW�pRW4PY5�PY6PY7PY84QO,�PFs�e1�� ?$VALU�3��̅4��0�Q�$��| n5	��C
1���0AN���R1�Rp�!��TOTA�LQ���7cPW�#I|�AMdREGENKj`b4�X!G�s�&��f�m�TRC�rKa_S���g``�3V'����c>�1E:3�@��ܚcV_H�@DA8}��`pS_YƱ�ڻ&Se�AR}�2��>@CONFIG_CSE��`RJ5_� ���Q�E� 4�{�O�v�k�F�PSܢ�F�f�C_YF��m���L�����(cMϰ���q�rd^⃁z��DEհ�2�KEEP_HNADD�q!��0�	CO�0+��A�r%�,�Of�
���q�,��1��,�REMC�@+����Bh����U4�e+�HPWD  �q��SBM!�D�uB� ,v�F1L�з���YN�p�M:�C���pQ�Er�� �l0DB�M�TRI�DA,�Bx� 0�K�TCLA�����U AYNSP��֡SEAꠁ�GK_P�Tn���B���RGIn�QSOL!UK ��P��)a&�$SC`0D�#ے�ALI�r���S�0�B#U�A}��P����� ���w1�q_�P�H�TIC�[�`�p[�REVIo��OLP���p��FK��_F�SSEGQ���b�*ց� c3�� �l0CP��T�U� MSEC��MN���̢�����`�R0�G����0O��1�$N�̡_�e�$�PA� j�P�vO�iP�MLr P�� ~�  �����e1���  $OW-����G����p� ��Hp2C�ĹAü�!ߤX�AX�Q��A7HI��6��ٔ@�2��Ϛ���BVF�EP���P�`�Q���H�ߢ�r��V�t��`a�B^"$4@:�Q������p�M���y�O��l""�SMH���<�M=�2� �@�L`UP_D�LY��ÆDELAk�>a2Yߔ��G��QSKI'�� i�P��O��NT\P�B��P�����`
� �P���a��v��l��� vP�ڃP�ڐP�ڝP��t�P��9���J2#�Z���yrEX@T�# z����z�.@�z��~� �RDCa>�� � ��0'TORq���	��!0�����SDRG��H���k���Gg��eE9R�qUBSPC�G�|z�?2TH2N�!�D�#�1� ����@��11�� �l�p2�F17��Ta��� Oѯ%��^������SD��VAHwOME�� �]�2e��k�}���������� ,]�3e�������0B �]�4e��ew����� �]�5e����*<W �]�6e��_�q���� �
]�7e���� //\$/6/ ]�8e��Y/k/}/�/�/�/ �p]�Sπf��  �AX^�u`� �]�ET��yp��m2.fk3I�O�p�:I0�� ��]�POW�� �� U0K���9x]�(d ���2�$DSаIGNA�L#gf�CJ�1@��RS232q5ӓ ����%8��I�CEt����³��I�Tq&aOPBIT�"cFLOWCpTRh003b��UXsCU+��M�SUXTđ��I���FAC1Dų%@ �T	@CHQ� �@{p�p��C�$��`�`OM,p_���E�Tޠ�sUPD�pA�3��p	@P�@�Q�W� !�(s�A�����)��.�ERIO�c��PT:p3T�2_`���Q/PDAMVWR����/9D��qV��6F�RIEND(�@�U�Fi��t�P���UMY�H�p@���GTH_7VTE�TIR���R��P�XUFIN�V_��ѥ�WA'ITI���WX���Y67fG27WG1��@�1SQbbgpp_�RE�O�_t��s�Q�`��[PC8�C�u��_TC3����p�e��GˀŲtqֱ@&Q/A�r�jQXp�EV��Ea����|���D�X s�ML����`��SX��(]E#T�CG3�WCPgw�s�|tD�LOCKkuvӮ�V��q�ta�$�f[���pkQe�RqY1}XlP2o[2�{3o[3}Z�y'�~Y�y�C�6.�s.�r$V�V��V8eVl���(�a�b!�غ��F�s ρ��fqB���`�R�4ɠ��E�$߂�S`�@a�Tu���PR�����uj�Sl�G��g T��D�� �����%s[��w���[��`�p�@|`�@��
��D�S�1� ؚ�R�_6�oQ���`RUMN��AXSA�`A�P�L�QV⮒THb��J���6�aqTF"�N|T���IF_CHeS���~�qU��6��G1@��0���� 6�7_JF?�PR�`����RTC� �μ�GROf�A�MB�Vq̐CrÃ��`UI�#���BU)cRSM0}��a`r�_W�P��TBC_P�PCMr��D��ЖLDR���ރoq��@��c�I�T�"��(���TA���� s���|� ��ҙ��� ���� �ݾ2�  2�� �S��g��	G| �Vд�}�I�8t�ˀ~�TOT��~��D젖�JOGLI�zC
`E_P��qBO���}����`�FK��_GMIR��Ѵ{`M>r&�AP]q��E)P�ҔJ�SYS�˂J�;PG'�BRK�bѕtߐ��I"1  N�pSY�x�D�A~��GBSO�}��0N��DUMMY15U��$SVVpDE_�OPoCSFSPDO_OVRU��� 3LD��óOR��� �NP��Fߑ�Ʈ�OV��SFڟ��.�F �́ճc8ؿQ˂�LCHDLz�REGCOV��[P��W�P1M��vձ�ROoC��r��_ ��� @��&`VER��$O�FS&`C;��SWD���r�����Rū�T�R�1W1FpE_FCDOƃ�Ӡ��B���BL�����1K0%�V@�Anr�@��b� �G�,�AM*Ã�D�Z��t�_M0�|B��3��OT$CA���DU���HBK�AЖ��IOoU��1qPPA�������������2��DVC_DB )c0�ё�21���́H��1P���H�3P���ATIOˀ�A{���qUtS젆6CAB�� nR�c7p���`S�oq���_�@ЖSUBCP	U�2��Scp�0�B��@sj�B��2��$HW_C_ dЧs�5�sAta���$U�NITb�\ U A�TTRI�i��C�YCLϳNECA�����FLTR_2_FI��8���6���Pǻ��_SCT6�cF_UF__��q
FS�1:�ZCH�A�Q�)9�qB(RSD���2x�ޣ�1�0;_TW�PRO���Ӗg@EM*0_��V�Tq� z���DIPҔRAIL�AC>��bMg�LOu��S��9�R܀��䁬����PR2�S�a��p!C$�$@	��F�UNC���RIN`�`Ԥ�'$fARA8 �b ��P#X0��P#gWAR/���BL�a�f'�$Az+v}(v(D�A`�Q!�(�#z%LD@�@��q�#��Z!ہ��#TI�5y����$�@RIA�A�2AF��P;A.3��45p�p�r@�MOI` ��DF_�P7��Ac��LM��FA�PHR;DYJTORG͢���fS� �5MULSEP�P����J���J������FAN_�ALMLVV�AW{RN	EHARDpP��E�Y"2$SHADOWl��/�?Bc֐@w@u�:�_m�ЖA�U�`�:�|@O_SBR&�E���JU &�|/!�CMPINF���k�D�!�CREG�pU��л�i�� �J��Q$;Q$Z�a�e�O�j��� ��EG�~���F*QAR�����2�q�7W� ,�AXE��R�OB��������R�_�]w�SY_�dQU��VS�WWRI�P=V5 �STR����T���E"W8�FT�qkB�`�B�P���V,�����O�TO�A8���AR�Y��3b���B�ƱFYI5�ܳ$��Kq1���Sa]�_�S��tEU3�zbXYZ'B:�j5�fOFF��Rb)zbnh7`B��"��d��V�  �cFI@� �gq��«�"���_J��6���y�$�a@dk6�qTB�)q�2arC� �DUt��DV7�TUR@!X
3�uAa�BX�P��IwFLg�Tд�7P�p�e�Z�û� 1�
8�K��MДDV�8���ORQy��V#�W3I��2�+�s0��h�à�Tz�OV	E����M� *��C�� S��
R��6@��*A�� W ��<�! �50���� �݀Q�*�������'�0S'���ER��Z!�	�E�PD��e�A����eH%t?g�!���!AX��6��!� �Ua���˙�1˙�` ʚ�`ʚZpʚ�pʚ��ʚ�ʚ1_�ʖ�0Ǚ �0י�0癮0���0� �0��0'��07��0G��d�X�DEBU-�$(!4C����vbA!B�����~�V��, 
#�Y�?�K�O W�#aW��aW��aW�Zq W��qW���W��:4fp�42���cLAB�b8I�) 6�GRO� Ir-L��B_�L��T ���`�@ �4�J�0�A<�AND���Z���e]�Ay� ���@~a`�ȳ!�ȡ ~`NT@~=!�SERVE��NP� $�pT Ae�!��PO��K@���-`�����_MRA�Q� d � T��e�ERRr2�00STY=�I��V�`���7�TOQ����LphP���RJ� ���|D@Q � p 84��Ԯ�_V1f���(�Ԥ��2��2����D@�p�H����$�W� ���q�VQ��@$���d0������OC�!P� � �COUN�T�Q  L�S�HELL_CFG�Q� 5!pB�_BASVCRSR��AB� ~SS�W�!h�1��%g�2���3��4��5��6ʋ�7��8��[�ROaO�0��Y`}`NLQ�lsAB�úi�AC-K4�IN�T� ���lpa@�0�_PUX�0@�OU�3Ps �l��I����TPFWD_KAR<�L�0�RE�Ę0PO`�! QUEr�t��� �r.@_AI@7�H��{`�D��EzbSEM�?Ox0)6�TYf*�SO��)�DI6��s ����b1_TM���'NRQg{`E�� (�$KEYSWITCH���I���HEupBEAT4�qE:PLE;�J�U��F���SN�DO_HOM20On<#REFe�PR�aP���Q�P7�C� O�1��v�O �;rK@0I�OCMgt��a� ��(G�HKQ� yDxat�RESUUB���M�"��w�wsFOcRCx�#\�G��OM;P � @��*3~@U�SP9P1��$9P3�4� yP�HDDNP�� �BLO�B  �p�SN�PX_ASP�� �0v�ADD�GA�$SIZVA$VqA:���0TIP��'#�A�� � $c�( �`bR�S��"QC7Л&FRIF���S����� NFjODBU��P���%�#�)��  ��i�P� x��S�IT�TE�sX��sSKGL#1Tab�p&���<3íP$0STMTd�qU3P&P�VBW���%4SHOW]5�AS�VDTU�� ��A00~Ħ2���7��7��7 �75��96�97�98�99�9A�9\P�7��7ӱ �6�`�7�C�3W�pH�9U1�91�91�91�9U1�91I1I1 IU1-I1:I1GI1TIU1aI1nI2�92�9 `@X�9�`@X�9Yp@XPI�p@X I2-I2:IU2GI2TI2aI2nI�^�h�93�93�93��93�93�93I3�I3 I3-I3:I3�GI3TI3aI3nI4��94�94�94�94��94�94�94I4�I4 I4-I4:I4�GI4TI4aI4nI5��95�95�95�95��95�95�95I5�I5 I5-I5:I5�GI5TI5aI5nI6��y6�96�96�96��96�96�96I6�I6 I6-I6:I6�GI6TI6aI6nI7��y7�97�97�97��97�97�97I7�I7 I7-I7:I7�'�7TI7aI7nD ��VP� UPDb���"+���
��0�GUN_C���s `�g�PUT'�cIN\�����AX�|�GO�U
GI~��IO_SCAw�ޒ0YSLOP�� � E%�"#��':' � d�� ʤ	�P��� �R��F��ID_YLj+�HI&�I����LE_g�V����$ ��SA���� hЂ�E_BL�CK��M1��D_CPU��F ��: &��Y�k�����b�R ;��
PW"���[ 	�LA�2S��h���RJ�FLO 5��5�đ 8�V��|V�Ĥ�TBC#��C!�X -$}�LEN��$}��D�RA��d!$��WI_��&�1}�C�2��AM�b��� 3�II�s ]���TOR���}��D����� LACEG��}������ _MA+ �J� �J�GTCVQ�r� �Ts sڒՈ����� �2��JF��$M�ԙ�J���0��� ���2/ ~0���ӱ�JK(�VK:�$�B�3,�J0O�>�J�JF�JJN�AAL�>�t�F�t�n�4o�5��N1�ܥ�d�N�ry�L��{� Tx��CF/!�T�v�M�?1�"B�NFLI�C�# REQUI;REEBUOy�n��$Tx�2�6��z� �x�. �3� �\rAPPR,�C���{�
��ENs�C�LOS� ��S_Mp� $ ���
�$���A?  �����  ����%���������s�VM_WRK �2 ��� 0  �5��)L �L	#�`������q���_���n�+5UX Ѡ;M_��� ���/B/T/7<I�)$ORk} �5/�/�?�/-?�;?1/r?�?g/y/�9DYN_�/�/�/e?O �/6O?O?]OkOa?�O��O�K��BSPOS�U� 1��� <�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
��8�B~�N�LMT������C  �1�I�N:�L�0�PRE_EXE]���l�.��AT}��J����LA�RMRECOV ���l��DLMD/G  "��LM_IF ��d�*�<�N�`��n��������ǯح�, 
�O���FNG?TOL  �K�@�A   4�F���PyP��N ?�������H�andlingT�ool �� 
�V8.20P/A�2E��x.p
�88150���8�0��334896�6��xis
991���pra�����rod7DE�3���pc 	}F�.014i��Y pFRL~�ld32����V�X��TI�V}�l�J�i�UT�O�� �h�P_CHGAPON=�З������L�1	� �������t�I��U� 1S  \����> j��4����VIQ�c߽�܇����� �3{���HG������HTTHKY �ߚ߬�����6�H�Z� l�~��������� ��� �2�D�V�h�z� ������
������ .@Rdv�� ����* <N`r���/ ���//&/8/J/ \/n/�/�/�/�/�/�/ �/
??"?4?F?X?j? |?�?�?�?�?�?�?O OO0OBOTOfOxO�O �O�O�O�O�O___ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ�lu*�TO�uχ�DO_CLEAN��|(��sNM  #��9�K�]�o�����_DSPDRYRL�'�HI���@(� ���%�7�I�[�m���������ǟ$�MA�XZ��t�q�q���X��t����i�PLU�GG���w�Å�PRUC��B�ϋޏ�П?�OD���(�SEGF��K������� '����%�7�o���LAP̏߮�Ӌ��� ����ӿ���	��-��?�Q�cϨ�TOTA�L�0���USENU̠�� �x���r�*�RG_STRI�NG 1��
��M��Se��
��_ITEM1�  ne��0�B� T�f�xߊߜ߮����� ������,�>�P�b��t�I/O S�IGNAL���Tryout M�ode�Inp���Simulat{ed�Out��OVERRɀ� = 100�In cycl����Prog A�bor�����S�tatus�	H�eartbeat��MH FauylD�M�AlerW� ��u�������������8�� �s�� �q�hz��� ����
.@�Rdv���.WOR�����X�/ /0/B/T/f/x/�/�/ �/�/�/�/�/??,?8>?P?b>PO��8� �0�q?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O_�2DEV�>,P�?_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso��o�o�oPALT D�a��o�o
. @Rdv���� �����*�<��oGRI���t��oN� ������ҏ����� ,�>�P�b�t������� ��Ο��b���RD� ���@�R�d�v����� ����Я�����*��<�N�`�r����PREG�n��0������ ��,�>�P�b�tφ� �Ϫϼ����������(ߊ��$ARG_��D ?	����k�� � 	$��	+[�]������^�SBN_CON?FIG kۊ����CII_SAVE  �������^�TCELLSE�TUP j�%  OME_IO�����%MOV_H8!�4�:�REP����X�UTOBACK��
��FRwA:\�� ��'`#������ ���x��15/12/03� 07:34:46���ت�B�T���x��숄����������"�����Pb t���5��� (:�^p� ���C�� //p$/6/H/'��  ���_��_\ATBC�KCTL.TMP DATE.D�l��/�/�/�/��INI��`��֞�MESSAG���!��s���|��1ODE_D&�����-(1O.P0> 4P�AUS�1!�k�� (7�:?��!�BPR;����@I>?�G=ԎQ���)�C��/��s9���? I�?>O  (On�(O :K$OZOHO~OlO�O�I�c4m0TSK  �s=���M�/OUPD�T'0�'dP5X�IS��UNT 1�k��� � 	� 
G ��` x�n��m ��"�����GP 7w�� TH� [ſ \q� M��G���b^�_�_GPX�N ��] ���Q ����?JT 7��_
� �O�_o o%oKo6ooo Zo�o~o�o�o�o�o�o �o5 YD}h �������� 
�C�.�@�y�d�����������P�)QMET�15]Pޏ7�ڏ [�F��j�������ٟ�ğ���!��E���S�CRDCFG 1}k���	�����@�����ȯ گ�����"���E�W� i�{�����
�ÿ.�� ����/�A�SϾ�Y���GR.PPQ?}�j kNAN�j�	��nz�_ED� 1t��� 
 �%-p EDT-k�b��ϼ߻�� @�-(����/����?�\�ϛ� ����2���a�EQPGPRE92�ߠ: 9۹�@$�k��ٳ�f��3\� ߩ���p;R<؅��� 7�I���m���4(��� ���d���Q�������9���5��d�A�� �������w��6�0T���T ��C���7�� � ��� /gy/����8X/��/�� ��/�/3/E/�/i/��!9$?�/q?�/���M?��?�/?�?5?��CR ���<ONO�O�O�?��?qO�?}���NO_�DEL�ϛ�GE_�UNUSE�ϙ�L�AL_OUT ���  gҜ�WD?_ABORT
_{��CPITR_RTN�  /����CPN�ONSTO��nT� ���$CE_�OPTIOkX��ƣPRIA_I�	PnU�P���PFFn�+[ڳ/��Q�_PARAMGPw 1+[�^�g�Qocouo4kC��  �n��`��`���`��`Ș`Ҙ`��`�`�`�  �D�`�`�`��`�d�`�m�a	���bD"p/�`;�pH�`Tpa�`m�pz�`�@ D��p�� D�`/�?���o>ogy��n|�`��`��`�� �C��p��p��p���p��`��`��`���`Ř`ʼpмp֪�pܼp�p�`� �����|;Mv� ���������1�� ŏ׏���I�[�m��� �������-�?�Q������	��i��PHE>�@ONFIGK_���G_PRI 1+[ �խ�دꯀ��� �2�D�V���K�PAUSPOS s1���S ,]E ������ƿ���Կ�  �
�D�.�T�z�dϞ�ЈϮ���j�O�Q��_�7�QO_MOR�GRP 2l }��0 B
�r�:� 	 :�R�@� v�dߚ߈�k������� ������2���h�V� ��z��:�L�������
�@�.��c�!݋���?o�o��`���0K���1r�����@�����������PP�½+U�` =Ua�-��k}��:
\�	�0P�N@f��5�Y`�53DB��+Y�I�2)cpmi�dbg[@m:o�  5�`5��U�ApG�k�`�$9��P	I�E�Z��`)  *�X�-/���0�0E�g/v/A/�`��fe/�/���/>?ud1:�/?��7"DEF ���7)�!c!b?uf.txt?e�?4 _L64FI�X ,  ��?�\�?�?�?�?&O OJO\O;O�O�OqO�O �O�O�O�O�O"_4_F_V~?MC�,P  d�_�_�UfS��t]��T�Ub=��fCpBp:�B��"�B��B����B�= B�a�C<z"�
�;�D�C���PD*��D#��ED)��Da��[�kE��E��=FhEF�q[F�=FH���	r�I���]���YF��T_�;�I���o�oM���o�lo~o�Y�oQ <u`�,� ����;���6g�� =<�	��U#����أ���ӣ�x,�;�C>�<����<�p  Dؾ�n��Dπ���fE�π�  E�ms�a�πz��C�  F�E��f�E��fL��  �>�33 ;���s�n,��@s�?5�@333�.��� A�UL��<#�
�2����/����~���Q���Q���E��� � H���1�9�J;#�H�2��Z��J�9�Q�e�w� ��������џ���B� �f�=���a�s����� ����ͯ����'� t�s�]��ρ��ϥ��� ɿۿ��5�#�v�2�RSMOFST c6>���9T1�P�DE !=�p�G���;�3�xU�O�>TEST02i��R7"r��|�| C4�ʀ���� ��!�C�BP���b� �aC�@i�-J:d�
-�I�_1�#7�-�T_�00PROG %�r�%v?��*�T_I�NUSER  ���(�C��KEY_�TBL  ��(����@0�	
�� �!"#$%&'(�)*+,-./0�12345678�9:;<=>?@�ABC00GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�������������������������������������������������������������������������������͓���������������������������������耇���������������������9�t���LCK���<��STAT`+��_AUTO_DO��%�INDT_7ENB� ���̟�T2�-�STsOP��SXCh�� 2$B� 
 8�
SONY X�C-56L輸�`߀@��ʹt( �АOHRC50K��o�7��Aff���// �>/P/+/t/�/ a/�/�/�/�/�/�/?�(??L?^?�TRL���LETE� ~�	T_POPU���-�T_QUIC�KMEN�4SC�RE�0B��kcsc�4��0��9��c_�4U�M�0U 1��_  <K�%k? gOK�EO�O�O/ÁO�O �O�DF<��_�O_P_��LStart �SM Comm �%IBSCMA�NS[_�NEnd�xV�@�U�0�_�]Us�er Cance�l�RUCANCA�C� o�L
�RRe�set�BURES oo3_E_�oYoko��o�o�o�o�o�@Z�ange�GZG_-A�_�ocuL ^��������)� ��_��ZVAG�_KONFIG.�RVW)��=�O�؏�s�-Dateie�L�%DATEI �1�����E��.�@� ��d�v�ß������П�"bMacro S�tep tt�PM�SK_}<��LW�ait Moni�tor3aSHTP �G�L�柫���������ZCYCLE �POW�PPWD������ DOW��%	#�_MAI�Nu�a�%Cb�NUA�L�?�ZCD���&��C�[�	���������?|(��$oDBCO� RI����5#DBLOVR�D�%�NUMLI�M��d���D�BPXWORK 1'���ϩϻ��������DBTB_N1 (7�P�Q����s�DB_AW�AY��GCP� ��=��3�_ALU��?3��Y�5���$�_DBG 1)ζ� ,I��K�!������
�͠벲����r�M� I�t�B�@��	�ONT�IM�7�����)��
)���MOT�NEND���RECORD 1/��� �����G�O�����"_��#v�������EXECU�TING

�� �	����)�P�������P�QELLED�������;������j�����������R d���s��0b�����  2���z/����Q_&�Vc�/�=������pj[� ��w��>/P/�t/_/��Z~
j�v�$�/�/�/�/c/?? ��E?��Q?u?�?�?? �?�?>?�?b?�/)O;O �?_OJO�?�OOO�O �OtO�O_�O7_�O�O m___,_�_$_�_H_����&
oo.o�_ Ro�_]o�_�o�o�o�o�?o�TOLERE�NC@�Bȉ�N�L����CSS_D�EVICE 10>�  üƹ Wi{����������sLS 11,}�K�]�o�����������rPARAM 2����Tu�TutRBT 2-4,|8��<I��� C�vd ����HR�&� & T�˴��?�g۶��p��  �\�  �g@��˴���A��F���p bR��Ɏ��?�B���vɅ�zɇă@��\�7�1���q@���Ɇc��Ɇ��� Z�l���������Ưد��7�� �m��C�wy�D�C�9���ѰA���A��ffAI��A;�33Ad  A�Ɍ��B�pѐ��U��̱C>��Bff�B���-��B*갉ֿ��ҿ��� }<� �b� K�@ S�D�ɍ )�K�]���E�sυϗ� �ϻ������>��'� 9�K�]�o߼ߓߥ��� ���������#�p�G� Y���3�������� ��*��N�9�r���_� ������������� 8!3�Wi� ������4 jAS�w�� �c�/�0/B/-/f/ Q/�/u/�/������/ ��/�/>??'?t?K? ]?o?�?�?�?�?�?�? (O�?O#O5OGOYO�O }O�O�O�O�O�O$_�/ H_3_l_W_�_�_�_�_ �_�_�/�O_2o�Oo -o?oQoco�o�o�o�o �o�o�o�od; M�q����� ���N�`��_��o� ����̏������&� o/�A�n�E�W���{� �����ß՟"���� X�/�A�S���w���֯ ���������T�+� =�����������Ͽ ��,��P�b�=�k� }��ρϓ��Ϸ����� �����^�5�Gߔ�k� }ߏߡ߳�������� H��1�C�U�g�y��� A������� ��D�/� h�S�����yϧ��� ������R); M_q���� ��%7�[ m����/}�&/ /J/5/G/�/k/�/�/��/��$DCS_�CFG 5�����!���dMC:\�� L%04d.C�SV�/�#=��A� K3CHS0z��/#>^?�?�  ����2�1�?�7� ��`iMU����(RC_OUT [6�%�!���/�!_FSI ?�I  �9#8AOSOeO�O�O�O �O�O�O�O�O__+_ =_f_a_s_�_�_�_�_ �_�_�_oo>o9oKo ]o�o�o�o�o�o�o�o �o#5^Yk }������� �6�1�C�U�~�y��� ��Ə��ӏ��	�� -�V�Q�c�u������� ������.�)�;� M�v�q���������˯ ݯ���%�N�I�[� m���������޿ٿ� ��&�!�3�E�n�i�{� �϶ϱ���������� �F�A�S�eߎ߉ߛ� ������������+� =�f�a�s����� ��������>�9�K� ]��������������� ��#5^Yk }������� 61CU~y� �����/	// -/V/Q/c/u/�/�/�/ �/�/�/�/?.?)?;? M?v?q?�?�?�?�?�? �?OOO%ONOIO[O mO�O�O�O�O�O�O�O �O&_!_3_E_n_i_{_ �_�_�_�_�_�_�_o oFoAoSoeo�o�o�o �o�o�o�o�o+ =fas���� �����>�9�K� ]���������Ώɏۏ ���#�5�^�Y�k� }�������ş���� �6�1�C�U�~�y��� ��Ư��ӯ��	�� -�V�Q�c�u������� ������.�)�;� M�v�qσϕϾϹ��� �����%�N�I�[��mߖߑߣ��$DC�S_C_FSO �?������ P  �ߣ�����"�4�]� X�j�|�������� �����5�0�B�T�}� x������������� ,UPbt� ������- (:Lup��� ���/ //$/M/ H/Z/l/�/�/�/�/�/ �/�/�/%? ?2?D?m? h?z?�?�?�?�?�?�? �?
OOEO@OROdO�O �O�O�O�O�O�O�O_�_*_��C_RPI����@_�_�_�_X_���|_�_o0o+o��S_GN 7��r`��2�[�0�1-AUG-24o 10:�`  ���{`3-DEZ-15 07:35�`�C`Ab Pj�,�i�a5n�`wa@�7����i�Z�X�_�o��VERSION jj�V3.3.2��lEFLOGIC� 18���  	Gh��Ny��]~�0rPROG_EN/B  5dEs�`�~sULSE  �cu�u0r_ACC�LIM�v���s��sWRSTJ3NT�wra���0q�MO�|�a�q/r�I?NIT 9=z����� �vOPT_�SL ?	;��
� 	R575�@ch�74m�6n�7n�50��1��#tNy���*wK�TO  �W��o�+vV"�DE�X�wdrbC`)�P�ATH AjjA�\KJBVTU�211160R0�1\ \  56S\ARG2\g�~m�KW\  Yt���mHCP_CLN�TID ?vEs� Go ǟ��I�AG_GRP 2m>���R�ؑ� 	 E�  wF,D�E(p ��D�5j�B�  �=�+�B�C�f�T�C�eEC�  C���CG�SCEZXB�Gm:j�f362 67�89012345����  � � A���A��=qA�A��33A�z�A���A��RA�A�ߠ����5j֠Ba@�  Aƌ`Ap��B�A�C�C��`B45l� 5eW�Ba
բ���{A�ߠ��ߠ�k����G��Aď\A��A�Q�7�� �2�P7�F�7�U��ߠχ�U�۠����������A�ffA�۠򠍿����ÿտ�[�_��Z�U�O��
AJߠD۠>*�8۠2�,O�&��8�J�\�V�`��A�[��Vk�P۠K
=AE�A?��8��A2��+ׁ
�Ϸ�������[��������x�q��j�c�\Q�;AT۠L��1�C� U�g�y�[���v�����Ѧ�-�=�G��I�>8Q�U�-�8���bq�7�Ŭ�}�-�@ʏ\����p����m@*�Ah��а��<�C�<��t�=�P=�hs=�ᗍP�-�;��
��<#��5lÐ�?+���C�  <(��U�b 4��̝�A����M�5iA@Ab?5����r� �����:��������5YkM	?Tz!�
�-��J�G�-�2��C`�-��xC���}�
���/G�{CEYA����ɦZH�����/��Ҧ��ED  E���D����m��/  8���T����D��𽲮 ?�~��k�f?��Ǹ�a��U�D�g�@ �à�"�`����o/��/J�/�"5iE)�0�	B���,��/?}/&??J?5?G?�?D`����ϧ�? �?�>�?OOD�V�� uWO�FO�O�O �rO �O�O�O�O_�O�O_ d_v_T_�_�_6_�_�_ �_o�_*o<o�_Ho"o �o�oto�o�oVoHO :%^I��� i����JT%�7 :��6�-��og�Iw� ����������	�� ��?�Q��ox������ ��ҟ�������>� )�b�M�_��������� �/��(�ϯL�7� p�[���������ȿ� ٿ���6�!�Zω?�? �?�ϴ��?�����+O =O/�Aߣoe�w��o�� ]߿��߯�����+� ��O�a�?���!�k� ��������'����� ]�o�M����/���g� ��G���$J5n �W����	�� "Q�CU7�y� ��Ϗ������ -//(f/Q/�/u/�/ �/�/�/�/�/�/,?? P?;?t?_?�?�?�?�? ���?O�?O:O%O^O IO�O�O�OqO�O�O�O �O_�O_H_wωϛ� �_�_���_�_��/ o/ooSoeo��9o�o �o�o�o�omoo�o+ =as�o�Y� �����'��K� ]�;������C/�_ޏ ɏ��&��J�y3� X���}��������� -��1�/U�g�y�� ����I�ӯ�ǯ	�� ŏB���f�Q���u��� �����Ͽ��,�� <�b�Mφ�qϪ��?�� ���ϙ���:�%�^��p߂�LU�$DIC�T_CONFIG� ?m�y�sVzPegWS�����STBF_�TTS  LT
�����VE�R��xQ����MAURST  LT��՜�MSW_CuF��@��ZP���OCVIEWf��A<������ ����������XR|� �#�5�G�Y�k���� ����������x� 1CUgy�� �����-? Qcu���� ��/�)/;/M/_/ q/�//�/�/�/�/�/l?��PM5�B<�xS��  ���;�SCH 2H<�
��yQSch�edule 1 >LW ��R�L�9ZP?�?M�HA8��1�?L[A�4>L�Ͳ2D�?�?�?O "O@OFOXOjO�O�O�O �O�O�O�O�O__0_ B_`_f_x_�_�_�_�_ �_�_�_o�TJafe�U4ueD5�9*o �9Dzhgno�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ�����5=`6�Je b�t���������Ο���	H�V��)�;�M� �?�?���?u�;oMoo ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ���_o �B�5�G��7�I�[� m�ߑߣߵ�����>� ���!�3�E�W�i�{� ��������:���� �/�A�S�e�w����� ��S��#5GYk }���I����92�?`�r�c��T ����ψ���� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?����?���� O(O:OLO^OpO�O�O �O�O�O�O�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o� &8J\n�� ���@R#�v� �?�?�?H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d��?�o���o�o�o ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L��o����� ����
��.�@������ 3. �� �6����v�(�:� L�^�p����������� ���� $6HZ l~������ � 2D��p�x �ߦ�d߶���� /"/4/F/X/k/|/�/ �/�/�/�/�/�/?? 0?B?T?g?x?�?�?�? �?�?�?�?OO,O�� P�O�O�O�O�O�O_  _f��b_t_�_���� �_��_z�V�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������PO8� tO�ODOv��������� Џ����+�<�N� `�r���������̟ޟ ���'�8�J�\�n� ��������ȯگ쯒O 0_b�t���������ο��F_�_"�4�F���4 ��_�_���_��:�L� ����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ^���4�F��V�h� z��������������� .@Rdv� ������ *<N`r��� ��R��B/T/f/x/ �/�/�/�/�H�?? &?�ϒ�c?��T?�,� ��?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ >���_/&/�o(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h� z���2/�/��&�8� J�\�n����/(?ԟ�`�5n�@?R?C�v? 4��_�_�_h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτ��_����ԏ� ������,�>�P�b� t߆ߘ߫߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�򏐟�� ��*<N`�� 蟢�� �2�V� ����ϖ�(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?�ϐ�x?���� ���?�?�?�?�?O"O 4OFOXOkO|O�O�O�O �O�O�O�O__0_B_ T_g_x_�_�_�_�_�_ �_�_oo,o��p�o �o�o�o�o�o � �bt� �6�� ���z?�?V?� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$��?Po X�to�oDo������̯ ޯ���&�8�K�\� n���������ȿڿ� ���"�4�G�X�j�|� �Ϡϲ���������� �o0�ߔߦ߸����� �� �F�B�T�f�� ������Z�l�6��� �������"�4�F�X� j�|������������� ��0BTfx ������~�0� T�f�$�Vhz� ������// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? r��BOTOfOxO�O�O �O�O&�h�__&_�z7����_��t_ ,��_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� �>�?�O&O�?6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ������2O�O"�4�F� X�j�|������O(_� ���`_r_Cϖ_4�� ��h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ���Я�����į�� ��,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZl�����/ /*/</N/`/ƿϢ/�/�/@Z8N_ �2�#? V�?�����H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_���_� ���_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L��p/ ԏ���
��.�@� �/�/������ ??� 6?ԟ�_�_v_��,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$Ͼ_p�Xϔ� ��d��ϨϺ������� ��&�8�K�\�n߀� �ߤ߶���������� "�4�G�X�j�|��� �������������P� �������������� @f���BTf�*9�/ ��ҟ����Z�l�6� ��0BTf x������� //,/>/P/b/t/�/ �/�/�/�/�/�/?~� 0�8?T�f�$�v?�?�? �?�?�?�?�?OO+O <ONO`OrO�O�O�O�O �O�O�O__'_8_J_ \_n_�_�_�_�_�_�_ �_r�boto�o�o�o �o�o�o&h"4F ����t:?L?? �������&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ^? o��4oFoo6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� ��Ro�o"�4�F�X�j� |ߎߠ�H������ �10��k \�្��ϟ���� �����"������j� 5�G�Y���}������� ������B1� Ugy������� ���Ͻ�!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?� ߻�OO1OCOUOgO yO�O�߻O�O�OYK� _o��R_��A_�_ e_w_�_�_�_�_�_*o �_ooro=oOoao�o �o�o�o�o�o�oJ '9�]��?�? �?�?�?����� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E��? �?�Oͯ߯���'��9�K��O{�����a���$DPM_SIM 2I���ʱt�������C&]Y&U� 6� 0� DϨ��q���RC_CFG� Jʵ�!�X�&]���ϸπ����� �5�6ᾰS�BL_FAULT� K��s�O�GP?MSK  &Tb����TDIAG �LʷհSQ���UD1: 67�89012345��xz޻P����� 1�C�U�g�y������������	��Y��۽@��RECP�ߪ�
��~�ܿ�ߴ� �������� 2D Vhz��������9�K�UMP_OPTION|�[��TR��}�_�1P�MES;J�UTY�_TEMP  ?È�3BȱЅ��A�oUNIT�|ׅ��YN_BR�K Mʹg�ED6ðZE|�'t�cԝx�TAT��EMGDI�[���NC#1Nʻ ���X/K/&^u�&[d ���/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O> COUOgOyO�I�!�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo�J<OFoXo jo|o�O�o�o�o�o�o �o0BTfx �������� �4o>�P�b�t��o�� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��,��H� Z�l���|�����Ưد ���� �2�D�V�h� z�������¿Կ��� 
�$�6�@�R�d�ϐ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������.�8� J�\�n�ϒ����� �������"�4�F�X� j�|������������� ��&�0BTf�� ������� ,>Pbt�� �����/(/ :/L/^/xj/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?/O2ODOVOp/ �/�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_O O *o<oNo`ozO�o�o�o �o�o�o�o&8 J\n����� ��foo"�4�F�X� ro|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�j�t����� ����ί����(� :�L�^�p��������� ʿܿ����$�6�H� b�X�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰������� � ��.�@���l�v�� ������������ *�<�N�`�r������� ��������
�&8 Jd�n����� ���"4FX j|������ //0/B/\f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�OO(O :OT/FOpO�O�O�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �?�_o o2oLO^Oho zo�o�o�o�o�o�o�o 
.@Rdv� �����_�_�� *�<�Vo`�r������� ��̏ޏ����&�8� J�\�n���������ȟ B�����"�4�N�X� j�|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�F�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ����� ��$�>�4� Z�l�~�������� ����� �2�D�V�h� z��������������� 
��H�Rdv� ������ *<N`r��� ������//&/@ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?��? �?OO8/BOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�?�_�_oo0O "oLo^opo�o�o�o�o �o�o�o $6H Zl~����_� ���(o:oD�V�h� z�������ԏ��� 
��.�@�R�d�v��� ����������� 2�<�N�`�r������� ��̯ޯ���&�8� J�\�n��������П ڿ����*�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮�ȿ������� "�,�>�P�b�t��� �����������(� :�L�^�p��������� ������ �6H Zl~����� �� 2DVh�z���� �$E�NETMODE �1O��  ����������RROR�_PROG %��%��:/G)%TA�BLE  ��%�/�/�/�'"SE�V_NUM �?  ��� �!_AUTO_ENB  %�$w_NO�! P����"  *�*20�20�20�20� �+10K?]?o?4HI�S�#���;_AL�M 1Q� �2��2<��+p?�?��?O"O4OFOt?_O�UT_PUT 2}R�=  @ٌ7����$_�"0  ��01��J�TC�P_VER !��!2/VO$EXTLOG_REQ�6s�9SSIZ_�TSTK;Y 5��RTOL  ���Dz�2�A T_BWD�@xP�&ܤQ-W_DI�Q S4�����VSTEP�_�_�>�POP_DO]_��FACTORY_�TUN�7d%iDR_GRP 1T�  d 	�O�|o�m`�[����N8��T&hB�( ����f�mc�o�mm`@���B$�Bs#���A�c�@9�xP�oB�B};�b�c��o�opG2k�h��Isy�A��et^s�p��k��?y��{r������ }/<`�>�q=�p����qs~
 G�y�q�uA�'�s��2_q{R }E�  wF,DG�E(pO��DE�4�D  E��o�D��w�m� }�C��N��B�ƹ��� ~UUU��U�U��0�B��� �E�@��� }OHcGP8��L�uS@�K�y�
 }?"�\���:G{:���9{�����Ԏ�l��s���ʀ���t��Jէpԏ�o�o00%U6�j 	��o0�ۏT�?�x�c� ������ү������ �>��;�t�#���9� ����ڿſ���"�� �X�C�|�gϠϋ��� ���������͟?�� ����%߇��߫��� �����,��P�b�M� ��q��Y���}���� ��:�%�^�I�[��� ��������� ��$ 6!ZE~-ߟQ� c�u�s�o D /hS����� ��
/��./@/��� v/a/�/�/�/�/�/�/ �/??<?'?`?r?]?��?�?�?�?�?\JFE�ATURE U��U�P	aH�andlingT�ool 'E al�lyEngl�ish Dict�ionary-A,� PaMul�ti Langu�age (GRM�N) t\ir�4D St@a�rd'F  pro�dAnalo�g I/OzG  �VLOA�Agle� ShiftzHl�.pc�@uto �Software� Update � \pk4�Cma�tic Back�up+Cirpk��Aground Edit @-A�@�uCamer�a�@F�I�@DPn?rRndIm�C)E��@Pommon� calib U�I S �@�@Con�QSPMonitoar,B�@�@kPtr%@?Reliab�@,B�ductDa�ta AcquiysoS,BAD p�P?iagnos�A�A�*D
PCV�Poc�ument Vi�ewe{R.@wc.��Qual Che�ck Safet�y[Q �Pl@Enh�anced Us��PFrP.@END�I5@xt. DI[O kPfi�T *`�F-bend`Er�rzPL�RdTKfgs�  ckToIcr��@3` BWD*DI�NT FCT�N Menu`v�S�AM@�`TP I�n�`fac�e{`t�\jG Pp �Mask Exc�`_@�EHT�`Pr?oxy Sv�T�A��QHigh-Sp�e`Ski;TdPc�s@�P7`mmun;ic�@ons.@�P\)qur�`�`�I.P��`�A�bconne�ct 2EWInc�r�`str�P�Vc�sgeKAREL Cmd.XG��e�sRun-Ti�$`Env�WK�`e�l +�@s�@S/�W-A�PLi�cense�S�Ve�tw�PZ`Book�(System)�*D   Q@AC�ROs,r/Ofgfse�@HTMH7`��@J��@ngQ@ec_hStop�atpp,�RPsiQ@iUb�K� p.f�@Mix�`�@�@'Gt`Q@o}d�@witchzH�93 R��pR�Q.�E� R808͆O'ptmڈPJ͆�`wfil�Vt I,`�τ�@gOw 0\t��PSB-T�`
SIP?CM fun�w�c�F OY�v�pRRe�gi�r=p�qGaP�ri�PF`� EL�SE���@Num �Sell�  oa�dx���"` Adj�u-p*DN@l@˕�J �\j76�tatau��Xx˕�Y  F`��`RDM Rob�ot>@scove�GA im�Rem4j�7anqG !b?�Servo7`��,B�!��SNPXs b�rzH596�`��CLibrFC۔H55��@ {����ԙ`��o�pt�`ss�agI� �aT�CP �C8�}K��/�I�m 1�p��MIwLIB!�.vrLP��`Firm�B'Gjq7á�`�bAccP2	U
��Q�TXJ��{55�Teln8�"�55 (��$A4��h�I)�`Torq}u�@imulayQ�Q tph�@Tou��Pa�q'GP��� P�Qփ&�`ev.�  i�USB� port SPi�PN`a�P P
�!1�nexcep���Y�n�S 9 R��i'G "L�`V�CWQr8r/rp�ڰ" ���P��\����@�ı���T��SP CSU�I��hc�P��XC���MA,`Web 3Pl�.�ER�`� y�O{�p̀/��`d�QLz`R�?�<ZC�@�e�GridD�play BAe���D�QJ�iR��.qJ����^��AAVM��IO`�pNa�PAxy`,B7�7����-ATXPL��+CHCSB9�-�2000iB/2�10 V b\��AOscii�aΒLŐp�P��L�c�UplŐ`'G���A���`opPBA 0���A�qW���ڸ�1�`CE�`rk�J�g R7PPR�UT����LQRT/�KeybowAMa�n^@v�:��PC�Pl� sd�by E-�c�Uol:@qQGuHwF|�C�P�@�@b�Q�kPss@tN@t�� Wtd\$�o�prE�ds@�f ��LQyc�@�r��ori`��P>�PCS Jo��sc`����@��a�Blu 4e��PH��<ZF�z,`D�@in N#ajy�.�5LPDy�܅�ifi�S 10i�@fDG@�p/��cUb�Outpu��B0�ࠃ`���im�iz��tm��KfA'xis7a�Q �����fm��s��  M�S��FRL�am�� ��P@HMI 7Dev�p (���� ␠P�aΐ��PM�h772�p.q/nn/C֐oޑ�@�J��x�o� �#1��u��773.�=��dЃZqRD��OD���Qb���C�o��qTXY�ROFI�NET�J "AM�0�d�Dp�GR�AM/JOG O�J����@ ! d�P�asswol�i�RL�`5!th����8�;SN�`Cli�Q#X�M ��SPEED OUTP���c`��� RHi��s=e8;01DpVAGn�rp��2"�!`vogi �7��BL$�#��3^.WGeavI�~*��V�~�64MB D p<Z� Ġk2FROs;w802DpArcҐ�viszS�*Aux<x�J&Cell�L6��9��OTsh�1(FM��@�<c݅]s�5�@pf�  m�7ty�@��@r2�@����(!9���� � p1`۔8I���w�./s��PR�� 2P��Q7�# e�@`�LR�ZvE% �Pu+DDf?�x�ʎPq`@5 fT1$G�T8���w40�  ���D�s��,���t�BOPT��pQ��SN`�`cu�[R�e� �p�Syn�.(RSS)$Ql�U�quiry`		 !0��?����� @8��t�
�QestSm0t-ESS�) ՠ�teHPWyS7@��miLjECSp�a_�N��h681�$r'�d�ib� LJ���P �cR��q��p�| iCA/l��a71{ap���=��!{aZ� EN9D  ��dpn����fd -�#V8.�x I�(��!EMZ$�EQ ñ�����LFREU J�e��d@a1 �#�s\0� + �� 8��when ar�g j�!���͡C-D�tip*=�Q�k�͡u8sd R.wSkif�WF,� oBCK TsAb��v!a�ung�pϠo��!r��P�!1��q68��I�Q�A �F�`b.Tig/�Td�(C� ix �up�� l�bof� GOسTo If��G�pQ�m�pOsfmn�p�s�t�Q� �:�-PS-�s�r�pL�@�Aff�.a.d S.PN�:FW-CHK �JG"�� ��\cdcCD:���SSTEP̢BW�D <�.Er.�af� 8xVa/g_C.l�j ��tsseJ�� Iss8`� iq�+P.A�lloc.Mem1.쀛k�29P���c I����w .K[��l Var.Sc;r &�O�����FB_CMB�lar��MNSࠏ�I��wr.�!FUNC�-Mx�R9`���	s� � S�˓k�n.�sMP 6��Z�c�md.er.-Pdl.�Prp��aEC�#rignǱ�& f�� }�TSHELL� Hebeat���No�.On�/��w.SRVOA ?!���,�9�m��� aw��6��Gu�nM.DO.@!.�Gen.�A R7�1l���?�.scr�n freeze� qP381�+Inv9`ig.���ch�peldp>Łx ABC&"g��p~�X '!.d��.�uP�p.��ar �gex.4�..abd PG�PX  R`�k�.��spddѐ4����p�� P}й�۳�3wp0տ��F�r���Rd�/�E�C�)��sg.E�;�!yaσ� Anl}���R788�ϻä0�W���������an#lg����`\	�+��Pp%�G�IS�A�cӈUr^��
Y�yߛ�8� J6�߷�(Li�n��S������o\aw�����ӿC��P9k=��ecoY�{��wmleu��MHy Dϳ�48 H��&��MH����Tِ���d "F�#�\mht�3�b�:�[��"AP�w�hto�t���B����ETU����ol$�.������l E=�5o�csQ�)��;���
4�54	5`�:�Ip�����H574��J�2���fa����`ą�j� ��ce�nl������H50��INT/��` -/�ķ�I/k#a�f/�z�55��-��/�#19��/'52�/�q0K��J?"MN�/�50��4�r~?�2�Z�!�?��u�4J�6_P�?�2��?t42�+D&0M%O;ūpBO� "@O��azO�B#ic���O�#0�/81�O�CpJ�O_']`��"_�Ӷ�8�ENY_lo�rϼ?-�_�1�O��R/��*��o#bx�Po��! ����- VUo��Rpoo8�ϯd2 J�o��Vi���A0�o�D�s_�.f ��ib���CLo/�_�2�O��Mp�;?�}v9m\cv��2Yt�T�T��Egnai��?]�����O�taX_N_4/a����a.@���cb_ -������e�;�a�9a���bsi��w���ޡ ���dӟ1ViAg|?�l/~/��r+��=���a�S�𯗟y
n�'�9�F���|�G�n�P��gί�ѿ  �ѐͿ�� A��53�1l~wO�O R�=ϫ�RS?�� F�6E09 ��W�o�0_P��dmTo¿H�Z�X/u� ��U�0����A���/��_��SEND���3� RX�r6��efJ9�Ϣ�AC4��P�_��mnm�~��.��x���CRL�*�\sIf�v61���j�/��6Y@i���fK�	�j`<��ߌ����ND����1p�f��fe(F<�?k�)�e�D�B/t�f���ZO�W q"H�O10F��ffe"L��5, �o�t\ha���}0���3Ttr��^�h6h�J�.z��ʕ
I%/���n�hm��buDE��?�ߓF ���V6��4Gc.$`j_��rl�� �/��0u?;��/�?YSC(?:?#F@f��_�e��9O+�H?�u74TO�D7 (� ?�����	�O^�L � feIn\/�gJ�5_�onO�VJ51��O*VI)�_�Dsf!m�_/E�_��e8�~_fxO48�O"ad$�2�I@/&�mn�o�c8� 4Z! j�o#csioF_X_59�?r3t8.o ingI 7�^p�o�t��|��5	P���!Lo�w(B��8O����PE��σ���}��o�Oȗ ����l_�/"/��a�� nit�/�Epld4_��!
�on|�8Ƈ��e G�JE�TX�:K���6c74=��߱N #`�n�gcr��/ߥ~u��ɯ{d.p����da���74�ﾯ`�r�0HG�q��2.p�vu�����/��\���_  :�2��7c.p�21k���3"�ݱR78�"�= P�0��J614��(�AT�UP  �OY�5S45��Y�6��s'��VCAM/�CRI<��=�CUIF��Y�s28O���NRE� t.vA���_ �`A��SCHO@��D�OCVO� -��D�CSU� p��J6�0^��0��EIOC6w�NT��54"�i��2��9�� Ski�SETw�q���1ûJ7��921@�M�ASK  K207PRXY�s��7�9�OCO{p�@1�3��ҵáQ�{pkmaY�Q�m�3�9�s���kckl�LCHN�=��OPLG�A�J�50~�r@I�HC1R�PE�I�CSj��`�l��Ђ�KAR��J{55^�rt FI�DSWo3�q����4q�f`nI�PRr����f����R��aU�CM���ӡP^�j�T��� f�9�1�v��L1�fи����v�209��P#RS*�́Y�9J�V��FRD����|�RM3CN���93R�n��|�SNBA�@1\�k��HLB��ME"��M��������q�m2R�in'�TCj�1�TMILC���A�2��p= )�PAб�vA�TX�Pkrc)�EL��Y��Ү�Y!Y�8E�rcfX�C�.���Y�95����95�f�f.v|�UECN���UFR����X��VCC��v \�VC�O��1.fL�VI�P.�735.��S�UIpL U��X�Ф�WEB�j��1�T��	���2n��g JT�CG���sIG��I�]% PGS�3% R�C.�I�s��\at.��H89v�8�Up1�X��@�H60.�LQ�l�R7�]�Rx���t�69���9������ "Cp�6Y1���J8��0FpЩ�v��q�7R�j6�70�3^�"FSEGY�8^��1��6~�J��HA�4��΀X��~�m�55v�ftp�$ J56������R�5��7%��R7n��tun0�98v����5e�U�82��sgt<�5���/�и��0.�70\$ R�55~�979��J�76R�O�0���5;73��J96ѱ����"��g��.�T"J0�6YF> ��4.�D)p� J���p�9������ ��57 �5@�A��~����\� ��^�b��]������в�Iß���V�5��tdf����^��Ĺ9ѵ�D06^�mch��"m�� ����wSVMr�men��LIr���v��C�MSF�V"� j���T�Y��6�I�CT�Oj�U����sgm2��5����NN��K0�f�mku8�ORS����%8R�$8��l�wEXT6 ��F\��I#OPI6 t� ����/�R6!!� ���PRQ  ��8L$���Sd2�w�2f��I�ETS6 U�SL]M*�svg�!6i��52^��� ��i�ase)�OA� L�)�RAN�&�3��sVA����IPN68H@.�=�EZE�0��  UPD~�%�U�M�C~�1�P1I�3E0}�3�@"��@~� ��@^���@�&�@��,��X�P1�
��B�.�9� �Bf��T20"�I#�@��al'��@����P2Q �B@��n�`�7P.��6Rn~�tol��P2}���P22v�#P2���m�sP&7P~�ks�e��sP�?�P24 ^�Fpl�7P^���P��v��S3U�kks��P27v�� ���P��0�B���P3����P4�1hk��P5�}�P5iQP5�I�a�P33��gkdf=e���������3J���U���sgk	t=e2 D=e�����!
=eI����k=e1" ������������ ��>��f5B��ABVe�� �e��e>���qB�e~A ��1����2���2��� �e��e����>eV! �e�A���B���ҶeJ!��tQ�f� �e2Q���=R�uJQ��hst. Ev�v ��m��e�!��ft�P�v�g�R�����������n����;4$��  =e"Z�<fak9�v5�o� orcm=e"C1C�U�܇cc�f�� �d9��f�����¶e]��g/`�:hm���hlo ����9�k
�T�֟螀}y����!0	�yfk�weyoY��ve����}���un<f�z���f�sub��c�fccce�+��fE�W�i�{�v��������Ğ�v����뛍iY�
!�s����� Di������f R�vT "�(�58��v� �vc�s/ "�:�� ag˗925"����f�26' �fr���E�^j�4ᨖ "DG�/�adg8v���on ��,vM�߄v1r��q�?dse��:�#di�����!�e�d -=ee	�yf��d�fN-��f82 vs�I�[�m�8v�Ϸe�l�Ϯ���sl8vG���T���ST��/�l �0�B��f�L���p�cdtHf����dg�߀b�����'�������d3ju8v{41�g�wZ��4�f51�v2�����n��ro�fst�K�nat�f0�� � �=e������PG`onSpox�, PȫNn�OFT|�bp�f�eqi�f��alu�f"WE��͌8vsweq��E�7`;tpȦu "p�&hV�n�wvK"�v��onf�vz��8ui��APF@�΀:�s��ftp�f����T������b�w8vI����&f4��-\��OT#/5-�dvG/Y/k'K93P�/�k9P�/�/� "K���/�  H55
P�!I1!IK946!I�!I=a!I�1!I�Q!I�3!IA!I9!!I�05!Iq�!Ii!�J �0!I9a!I�0PJ�!IaqJ"SC!IY11J�!IP� !Iua�J� !I�qZ�!I���Z��!Iin.@J�_we �_�_%V��1_X�p�_��Yu�J]_o[=o?[ld_o�[_Ko�_�_#G�homj)�!Ig\ff!IU�1O#G��O#Gaxtd�O�O�o0�oa��o�Yax�o�'��4ASysw�as���#�F�ztp�J}1Q�h��FGMQOcG� �J-^;h5 ZAR"�k�0�!Inrg�j-M5110�O_ė " �-�0\s`zyaJ��J�MNI��Hfmn���)1Z]���NJP9"q�cGmnm�Z�Mb^�0�~_�[t ��@�1���qOÏEWT0Z`�m�������PD ��]Mpsy����dFFί�Zrl��0��0�FRA��`zm��2* E����er�ZM�&_�RSo�1�y���� ��Ɵc� ��?K���CLPZ�}tps8Z]�o�PMA���Ims�J����n���ym���#�5�7�Y��8��}��GRD��]B��bd!�-R"�]��"�DN0!��"�odt`�-B"�-�"�=�r�P"�r^�"�-�"��� "���"����S��"���r"�n�i1�C��E9M_�!�emd�������������� �
ssp
t Iy)q"�asde!�w !  � us@
�rsal!�!
�IAR831di�n$�m� P�ar��b�\sr�g�F  !�
�! s�ServޡIF O�37{ R�Load�7rvo�I)o��R�def.�s�+! mi*G C���0*8- !+��ޢng M�E,� P���A�gc�o��pL�migp*~F�*� ��q�=0�f.s*-���0e�NDO;fdv�+ -�+ive�ܝ²)691!:RI�N�701�pti*��2I} �+�j`:j703�* �OpJ�?O!K3�set,!?�O�?��+�M� �:dnp*ER{ J�1 R6Z�T_+ (MI�voi@* "�+��?�$H6�*g.f@*Jwog�R52��che@*^  j�r��_Wog�*lin=k�k I/Q_#H� J5A;P0* J8�j/O,���B);cl�*v
�J~`ހ*pprx�Jrox0z�o�k J68o ��B(�P :]�r/�(�mPj��Simp��te�+R609¡[L�z��o�ZtorPjspa*tch�J�th *AST kH�ST�*794�zi�n�T��a?Sta^ *�Aϋ`���b��_�5p.pJ�CP�|58�J�M�odbAOSObt8�;��+PRO [ �O"�930�;�/:�30\0�_�+FS�W�}�o�h9pZaqm����*t\j�hp J�? ��Co/�]]=-ol/�N���=�8\gpJ�0���R	Co��e�Np�}_i0*VM���_�[�0� j92o��P�ceaN�:�M~P0:(N?+� WC�O�)dnw��EN�:��- �L�I/F kJ5���r w�:ar ��rj?�}@�;cm�n a0�M=�.�0����U�g�)�c��p* j6�TorP_R�D)��=oOkM�oCR HA� H�j�=1\�;�=�@�*^�@*h f�z-@��o82 (a*r : �����������P:982�*0�0�B�
�'0_�Sq�����������0��P:580��*1�\ pa���j����5����W!e�mOkm�4�\n�9-A���804 j΀& �usO�-�\�ڍ�a*n p:�M���ZJ9ϫiM !
mq��M`q�p�zj~,mo�o� �����@��i7 �J�� zm�/cυ(� l6�
H5;80Y6 �M�54_�nN��`�cz\P���  STD��?LANGK0-��1Em�C%E��%E67�1%Em�%E (S]emFCha%Et��%E�� %Ej]@%EM��%E��6IG!�F- �wO)A-%ECmp%EJx�HM�%Eg SV%E�o H�F>�PIGPHF�!%Eh�p�H�F��8�Fn�mFfunIO��83`OrCt%Ect�io�F=0%Em�%E8�3\s%Eq�G83��H8�FD j%Eu�tpumF] �G19BUF9/@"U=�%E(`�!V%`mF��%E�@pf8�46\%Em�mFj8y4%Gg M90%EHiOpg2hm!%E��%E00iA%Ept�,�F�%E͑%Em94l%E��f>��fZ_�l_~XInt�FQI7�58�_
�FXfrfqaPV�_'C58\Tv�k75�o��FL-��O;�-��o�k-ne|�V=1RBT
9r�P_�9\f0p_���S_��p9OP�TN�B5��Saf=e��by F��QBN��586<@��6q ��=љ����э�]���������!���r4���]r��ir��}R�� �Tri�����25 H��PRA����Io�Q��r6Q~�C��NQ��gRq��]!���q����O��!A�� ���F�Q��j62��!w ma��- P��gnapȆ��96�iBZ�(;����/�%�DPN)@ �е�I�8��U���Plu������B��7҂��݃ۤa���1����������p@Β���Ҭ�P�IZ��]���������R75�4�k�I�0�bsk@l�����]�萷�1^����sr�ts/A��Dp]�妕���J91��8�!ƺ�CUSa���g�itpl�g��gÜ��g�sdm�g�S�ys<@gþ��R {SMe�J737��0Qf�P��DsK�g����Ie���e�\sy�(���s���menqueŎ���Dat0��g�etw��Ň�7�40��i�g� (D�T�.bO���Par e�9rf�Er��Βg�=��g�I�s�n�s� U1pe�m�g�07{��ԗR72m�9ǁg�4� R8��7�pR"<m�E�7 (AE�j�I,E�>0
E�f�dE��in\P��RRas�cbE��BR- T�OE�rts�%�R�R�D�R617E�01싰j�R6��609���1�j�TQS]�f�o`R�BR�B6�qsx4���U�! cnE�OContE�prE�<m�R56 JE啲�RJ756E�lNO�Rc5PE�q��"q.��nsvE�E� 5��� E�bdr thƓ�iv��ْ��55����0����58��J̋��88��"OB��bO穒�淐^�NQ&B$mb����v�B$/h848E�2�a��� 48s�UbB&���9 E�H612�E�w� (��250�F]Y�j�f�
\sĈ��N��i�h6�1��200��RS H����L�3��B/1ybB$�b��\]�b��ae�G�K� I/��E	79p�P�$iBj�(EG]�e��/$*gd\glY�#�gd�cy�� C�'Tr�p �22�煒�4���4y;clX&ack8�/?5t8&�$����U��er|����4��H��CVT��KL�� PH(���L���6`90�30�8>�&^94ǀ^M�����:E3 �  �]$CL\�����9��$]Z<q@]9M �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿���99G�����$FEAT_D?EMO U�@�A��;�   �N�D�Vσ�zό� �ϰ����������� I�@�R��v߈ߵ߬� ����������E�<� N�{�r������� ����
��A�8�J�w� n��������������� =4Fsj| ������ 90Bofx�� �����/5/,/ >/k/b/t/�/�/�/�/ �/�/�/?1?(?:?g? ^?p?�?�?�?�?�?�? �? O-O$O6OcOZOlO �O�O�O�O�O�O�O�O )_ _2___V_h_�_�_ �_�_�_�_�_�_%oo .o[oRodo�o�o�o�o �o�o�o�o!*W N`������ ����&�S�J�\� ����������ȏ�� ��"�O�F�X���|� ������ğޟ��� �K�B�T���x����� ����گ����G� >�P�}�t��������� ֿ����C�:�L� y�pςϯϦϸ����� 	� ��?�6�H�u�l� ~߫ߢߴ�������� �;�2�D�q�h�z�� ����������
�7� .�@�m�d�v������� ��������3*< i`r����� ��/&8e\ n������� �+/"/4/a/X/j/�/ �/�/�/�/�/�/�/'? ?0?]?T?f?�?�?�? �?�?�?�?�?#OO,O YOPObO�O�O�O�O�O �O�O�O__(_U_L_ ^_�_�_�_�_�_�_�_ �_oo$oQoHoZo�o ~o�o�o�o�o�o�o  MDV�z� ������
�� I�@�R��v������� ُЏ����E�<� N�{�r�������՟̟ ޟ���A�8�J�w� n�������ѯȯگ� ���=�4�F�s�j�|� ����ͿĿֿ���� 9�0�B�o�f�xϒϜ� �����������5�,� >�k�b�tߎߘ��߼� �������1�(�:�g� ^�p���������� �� �-�$�6�c�Z�l� ���������������� ) 2_Vh�� ������% .[Rd~��� ����!//*/W/ N/`/z/�/�/�/�/�/ �/�/??&?S?J?\? v?�?�?�?�?�?�?�? OO"OOOFOXOrO|O �O�O�O�O�O�O__ _K_B_T_n_x_�_�_ �_�_�_�_oooGo >oPojoto�o�o�o�o �o�oC:L fp������ 	� ��?�6�H�b�l� ������ϏƏ؏��� �;�2�D�^�h����� ��˟ԟ���
�7� .�@�Z�d�������ǯ ��Я�����3�*�<� V�`�������ÿ��̿ ����/�&�8�R�\� �πϒϿ϶������� ��+�"�4�N�X߅�|� �߻߲���������'� �0�J�T��x��� ����������#��,� F�P�}�t��������� ������(BL yp������ �$>Hul ~������/ / /:/D/q/h/z/�/ �/�/�/�/�/?
?? 6?@?m?d?v?�?�?�?��?�?�?OO2M  )HHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ���&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ�����>0�  1�,� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r����������̿޿���&�7�:�-�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� ������ *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t��� �����������(� :�L�^�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8I��$FEAT_D�EMOIN  V:D�h@�3@PD_INDEX]KlA��P@ILECOM�P V�����AkBKE�@S�ETUP2 W��E�B�  �N �A�C_AP2�BCK 1X�I�  �)MA�KRO900.T1P:G_3@%�E_B?Z&_c_:G�E1__UT1]_C_�_�_y\2�_�_UT2�_�_1oDnoy\3ooUT3eo Ko�o�oyU9H�lJ3@�@8u� (��^���)� �M��q������6� ˏZ�ď���%���6� [��������D�ٟ h������3�W�� P������@�¯�v� ���/�A�Яe����� ��*���N��r�ܿ� ��=�̿N�s�ϗ�&� ����\��π��'߶� K���o���hߥ�4��� X����ߎ�#��G�Y� ��}����B���f�@�����1��K�@P�O� 2�@*.V1R:���RP*����`#S����yUn�PC��<RQFR6:��4��X��T|@|��y�_@I�xVG*.Fq�%Q	��<�`�STM ���" ���RPiPend�ant Pane	l��H�/�/p�Pi/�
GIFs/��/��/F/X/�/�
JPG�/!?�?�/�/�q?��JS{?�?RP�73�?O?%
JavaScript�?�/CS�?(O�O�?� %Casca�ding Sty�le Sheet�sTO~P
ARGN?AME.DT�O�l�\�OUO�1�D�O��O	PANEL1�O2_%�_[_��_2P_�_EW�_a_s_oZ3�_:oEW(o�_�_�oZ4Xo�oEW�oio{o�DSH�ELLp�A %�+rCm���GZG_MENUE0�-O�u�q���EE�INGAB�J�%�3�K�L�����vS�UMM_VAG.ID>?�O:���������yTPE_STAT:��;�S�y������E;�INS.X�M[ҏ�@���o�aC�ustom To�olbar ��yPASSWORD�o~U�FRS:\C��� %Pass�word Con�fig���G�CONF1��]��Aǯ�����,��yEXTSERVOC�U�K�c��������UIO_S3ET|��%�AϿ�	���4ϣyVWEMZROUS�e�S�kϰ���ϼ�K�AGV�UP[�m����ϙ��@� ��d�߈ߚ����M� ���߃���<�N��� r���%����[��� ��&���J���n��� ���3�����i����� "��/X��|� �A�e��0 �Tf���= ��s/�,/>/� b/��/�/'/�/K/�/ �/�/?�/:?�/G?p? �/�?#?�?�?Y?�?}? O$O�?HO�?lO~OO �O1O�OUO�O�O�O _ �OD_V_�Oz_	_�_�_ ?_�_c_�_
o�_.o�_ Ro�__o�oo�o;o�o �oqo�o*<�o` �o��%�I�m ���8��\�n�� ��!���ȏW��{���"��$FILE_�D�� 1X������� ( �)
SU�MMARY.DG�#��MD:W����s�Diag S?ummary����=
��SLOG��p�Ђ�۟�����so�le lo����T�PACCN�v�%�^�����TP A�ccountin�=���FR6:I�PKDMP.ZI�
�j�
� �����E�xception�$�ի��MEMCH�ECK���������/�Memory �Data����� �)��HAD�OW������)ϸ��Shadow C?hanges,�ߴ��O�)	FTP����χϲ�1�m�ment TBD���ܷ\+�)ETHERNET���͎f���3ߪ�Ethernet 3�?figuraC���~��DCSVRF��p�Ϝϵ߸�%z�� verify �all��cĐe�u�DIFF�ߓߥ��:ﹰ%��di�ff<���f�z�CH�GD11��*��c Q�����9�}��2����C� 8��j���GD39� �2��� Y���}��UPDATES�. ��ЋFRS�:\L7�Up�dates Li�stL͛PSRB?WLD.CM{ό�7�N0�PS_ROBOWEL��g�:SMp�)��M���/Emai�l��aïcį ���Տ���� /�� $/�H/Z/�~//�/ �/C/�/g/�/?�/2? �/V?�/c?�??�??? �?�?u?
O�?.O@O�? dO�?�O�O)O�OMO�O qO�O_�O<_�O`_r_ _�_%_�_�_[_�__ o&o�_Jo�_no�_{o �o3o�oWo�o�o�o" �oFX�o|�� A�e���0�� T��x������=�ҏ �s����,�>�͏b� 񏆟�����K���o� ����:�ɟ^�p��� ��#���ʯY��}�� ���H�ׯl������� 1�ƿU������ ϯ� D�V��z�	Ϟ�-ϫ� ��c��χ��.߽�R� ��v߈�߬�;������$FILE_7 {PRF ����������MDONLY 1�X�� 
 �q�H��l��y�� k���U������ ��� D�V���z�	�����?� ��c�����.��R ��v��;�� q�*<�`� ���I�m/ /�8/�\/n/��/ !/�/�/W/�/{/?�/�?F?��VISBC�K#��2�*.V�DM?�?0FR:�\f0ION\DA�TA\�?)20�Vision V?D file�?�/ OO3?AO+?eO�?vO �O*O�ONO�O�O�O_ �O=_�O�Os__�_�_ d_�_\_�_�_o'o�_ Ko�_oo�oo�o4o�o Xojo�o�o#5�oY �o}��B�f ���1��U��������MR2_GR�P 1Y���C4  B�r�	� .�ҏ�πE�� E�@��������πOHcGP{&�L�uS.�/K�y
�?�J����π:G:�r�9�{��~��A� � ����BH̃C�{�NƕB�ƈҕ�΄���π@UUU�UU��S��΁>t�>S���=�h=����>�=���;b��B:{e�g:�sX:+�N:I9���2���V����̃E��  F,D�E�(p�D����0E;��5�D��=��< Əd������������ �οϊ���:���_� ��nπϹϤ����� ���%��5�[�F�� jߣߎ���J�\��߀� !��E�0�U�{�f�� "���F��������� A�,�e�P�u������� ��������+( a�߂�d��� ��'������ ������� �#//G/2/k/V/h/��/�/�/�/�/��_C�FG Z��T ��/5?G?Y?��N�O ���F17469w ��-RM_CHKT_YP  0�r�h��00��1OM�0�_MIN�0r�����0��X��SS�B3[�� �
De; C�)O8K��TP_D�EF_OW  �m���PGIRCO�M�0aO��UNC_�SETUP  ���%O�O�O�O��G�ENOVRD_D�O�6}�mEUTH�R�6 dUdT_�ENB�O PRWAVC��\�7�0 ���_�/�_�_p|O�_� �_ (o�_Lo^o�_mooo �oyo�o�o�o�o$�o HZ�o~��3y�dQO�@1b���r��eB�8��^���
��F� � ��à?ϝ_�D��Zr�t �>0��x��g�f��B���r�	�y���!�&���"�D�F�x��������Z� Ԇ鏓���}1\�>� �:�\�^�����˯Ɵ@����ܯ ��At� V�'�R�t�v���ѿ��ޯ����OGRSMTkScrY�p�0w��m�x��$HOST�C21d�y�0�IQa}U@k����q��k1�72.26.18o.230��e�� *�<�N�`�n�e�ϒ��߶������� e	�cfg_fanuc���.�@�R�b�� Eu���eB���إ�� ������(�s�L�^��p�������9�	anonymous�� ����e�w��� t�������� =�(:L^��� �������9K ]6/qZ/�~/�/�/ �/q/�/�/? ?C/ D?�h?z?�?�?�?� //1/3?Og/@ORO dOvO�O�/�O�O�O�O �OOQ?_<_N_`_r_ �?�?�?�?�__)Oo o&o8oJo�Ono�o�o �o�o�__%_�o" 4F�_�_�_��o� �_�����o�B� T�f�x�����o��ҏ ����Sew��� t��������Ο��+� ��(�:�L�o���f��������ʯ?Ώ�EN�T 1e��� � P!a����� 	�F�5�j�-���Q��� u�������Ͽ0�� T��x�;Ϝ�_�q��� ���Ϲ����>��� t�7ߘ�[߼���ߣ� ����:���^�!�� E��i����� ��� $���H��l�/�A����e���������QU�ICC0����!�172.26.1O8.851G#���	2�s���!ROUTER��!7`��?PCJOG7�!192.168.0.10~CAMPRT��c5 x1���R�T ��%/�NA�ME !��!�KJBVTU21�1160R01R�S--KU1�S_CFG 1d��� �A�uto-star�ted2�FTP=��!T�V��/��? ?1?C?U?��y?�?�? �?�/�?f?�?	OO-O ?O��/�/�/�O�?�/ �O�O�O __�?6_H_ Z_l_~_�O#_�_�_�_��_�_o�o 	SM<����O�_to�O �o�o�o�o�o�_ (:Loo�o�������� �2�D� �ZC��og�y����� ��Z�ӏ���	�,�-� ��Q�c�u�����THC� ���'�I��4�F� X�j�5�������į֯ ��{���0�B�T�f� ��ß՟��ҿ��� ��,�>�	�b�tφ� �ϻ���O������� (�s��������ϔ�߿ �������� ���$�6� H�Z�l������� ����5ߛ�Y�k�D�� ��[������������� ��
.Q���dv�����4(_ER�R fF*��P�DUSIZ  j\ ^w���>?WRD ?�%:���  b�ackup�guest�Tf�x��3&SCDMNGRP 2g�%w� �:��\ kD?K� 	�P01.05 8��  ��  �� ��]  �Nw��� ����y���2; �����������+-(� g ��v@<+/�=&9���V����? �S/�  
�  �s#�� �{/�j���(���S�#+�� U�/� 5�n 9S`��d�/!/�/E/2���1234567& �?��?�?�?O�?*O ONO9O^O�OoO�O#; �O�O�O�Oy?�?�?F_ �OV_|_g_�_�_�_�_ �_�_o�_	oBo�Ofo %o�o__)_;_�o{o �o,)bM� q���Io���|(��_GROU�Uh�	-0�	��!1�cz���B�QGUPD?06��C�V��TYv �� �TTP_AUTH� 1i� <!�iPendan������!K?AREL:*$�-�?�KCT�d�v�L��VISION �SETM�ԟ��\ J��ٟ�I�'��?� 9���]�o��������CTRL j����
 (PFFF9E3ȯ�8�FRS:DE�FAULT2��FANUC We�b Server2�
�,>۬�����Ŀֿ����WR_�CONFIG �k� f2��I�BGN_CFG �l��2\ @�\ <#�
~�BH2|�C��?4:�~�L�DEV�`��|V�� IO ma��I�EXDAT �n����EXFLG����T�FIL �o����O�TP �pYݮaR!B���R ����	MERC�ATOR!REC�O�� "R_ACH�S��ISTW*��V�,�V� "SEN{SP��TXQ��990 	Keine 0�k� h�\%IB�SC����M�4�8�2@�EW�𛩀�TĿLMTN  ���� ����������l�X�SBAD��� 7�^�x�T�DL_CPU_kPCQ�\B�B���� @��[�M�INd� =��-T�GN��O�H����рINPT_S_IM_DO������TPMODNT�OL�� ��_PR�TY����Q�OLN/K 1q�@9�K]o���M�ASTE����SLAVE r����OZ���UOxv �CYCLu��$�K�_ASG ;1sY� �����a�՗�~���`�$0c�������a �������%/0/ B/T/f/x/�/�/�/�/ �/�/�/??,?>?P?�b?t?�?�XNUM���扜�O_IPC�H?��O_RTRY_CNQ�I�D�QN؁��8�� �Z�t��FO��T�SDT��OLC�������$J2�3_DSP_EN�B�0�ь@OBP�ROC�C���	JO�GI�1ukL�ad8�?����O��??�ۯ4_�pQ J_o_�_�_R_�_�_�_d�_�zO�y8!�O -oo)_;_�_�o�o�o �o�o�o&oJ�B1+oeNaoso�o �����(�:�L�^�9���BAc���� �����*�<��� `�r�����q����C��8��?�BPOSF�O~F�KANJI_� �K���RE_�.Av�/��/�����KC�L_L��2�?�EYLOGGIN7��М����$�LANGUAGE� ����EN?GLISH ١��LG-Bw �S���*S�x ����B�����S�'� ����Z�MC:\RSCH\00\X������ISP x���؊�⍊�ߡOCl���Dz���Aݣ�OGBOOK 	yYݟ$�챟Xx�	��!�]�x����`͛ѧ��ه	ε��>��ϼ̲�_BUFF 1z(�ϟ��ߞ /��K�]ߊ߁ߓ� �߷���������,�#� 5�G�Y��}����ǿDCS |ؽ =��͑�L����$�6�H�Z���IO �1}cJO����� �������������� #3EWk{�� �����/�Cn�ER_ITMhNd������� �//,/>/P/b/t/ �/�/�/�/�/�/�/?���qSEV@�.mTYPhN�l?0~?�?=��RS�0��|��BFL 1~|�@��OO(O:O0LO^OpO�?TP��y�[2��NGNA�M]��6ˢ��UPS�c�GI�0c�����A_LOADPR�OG %�%�UP051}O��MAXUALRM�,ܑ��筥
DR�A'_PR�Dܐ³ڑDPCf�ع�ͪ_�$�;Y�P_GRP �2��[ �S�2�S�	[1�ڐ+  ��_���R#oo  oYoK�Go�oso�o�o �o�o�o�o*< `K�gy��� ����8�#�\�?� Q���}�����ڏ�Ϗ ���4��)�j�U��� y���ğ���ӟ�� �B�-�f�Q������ �����ǯٯ��>� )�b�t�W��������� ���ݿ��:�L�/��p�[ϔ�=WD_LDXDISA�@+;l�MEMO_AP�@�E ?�K
 T������&�8��J�\�n�DPISC 1��M��ϻ��T�Q ���߅����2��V� h���w�K������� ��
������R�d�O� ��o���-����������*��C_MST�R �,=ISC/D 1��͠� ����� :%^I�m�� ��� /�$//H/ 3/l/W/i/�/�/�/�/ �/�/?�/?D?/?h? S?�?w?�?�?�?�?�? 
O�?.OORO=OvOaO �O�O�O�O�O�O�O_ _<_'_9_r_]_�_�_ �_�_�_�_�_o�_8o�#o\oGo�oko�o:MKCFG �X��ogLTARMu_�b�X�b �c�� (t�b�_GRP_DO ��X�a���?�L��uq�>k�����o$?MMETPU��Xs���`	NDSP_CMNT��`�Q  �I��q�al�|v��POSCF"�9�f��RPM!���STOL 1�X� 4@�`<#�
���a�� ���� �"�d�F�X���|��� П��ğ����<���0�r�\��SING_CHK  %��$MODAQ�c���o>�i��DEV� 	X
	MC�:C��HSIZE��͚`Ȭ�TASK� %X
%$12�3456789 �M�_���TRIG +1���lX%�ܪ� �c��Կ����˿Ͽ� <����7τ�+Ϩϋ� aϣ��ϗ������/��YP���`��E�M_INF 1��w `�)AT&FV0�E0%ߜ�)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ������H�� ���D���AL�t� /������ ���� �߸�����M� �q��� ����Z��������� %����[� �2�� ��h������3 �W>{�@�d v��/�//f@/ e/�/D/�/�/�/�/ ��?���a?s? &/�?�/�?v?�/�?�? O�?9OKO�/oO"?4? F?X?�O|?�O�O6O#_ �?G__X_}_d_�_�n�ONITOR=�G� ?��   	?EXEC1�c�RU2�X3�X4�X5�XTp��V7�X8�X9�c�RkBOd�ROd�ROd bOdbOdbOd%bOd@1bOd=bOdIbOc2VhU2bh2nh2zh2�hU2�h2�h2�h2�hU2�h3Vh3bh3�R���R_GRP_S�V 1�q� (�d�:2�?�BM��;���@I�7?�=ԍ9�Ze�C��c���z�����U7�_�D@R���PL_N�AME !>��Y��!Defa�ult Pers�onality �(from FD�) �TRR2hq �1�����Y�  	 d���ŏ׏��� ��1�C�U�g�y��� ������ӟ���	��+�2��K�]�o�����@����ɯۯ��<:� �)�;�M�_�q�����৿��˿ݿ�  � �\  ��  ��  ���  A�  BU�T���
���
��@��  �Y���B�p�o�  C�C��P Dz  E�;� E@ D��c�C�J�q�X� �d�Y�p�t�l�`�u��e���È�d�\�]�E�/~ĉ�\�����`�@o�e��`ż� �E	נŌ��^Ì���t�\�@�T�|���EZ���å�]�|�Yũь� EY��ߧө���`���¡���]�����0�������� /�� ������D�M�a����q�]������T�E� ������]� �/���-�O�Y�M�s� ��������������� V�%ثD��E��x �  �s�>P
�d�tl~c���! ����� 6 �'EK i�������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? -�F?X?j?|?�?�?�? �?�?�?�?�O0OBO TOfOxO�O�O�O�O�O�O�M���O\)� _E_���c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�oR_�o�o �o�o�o%7I [m�����o ���!�3�E�W�i� {�������ÏՏ��� ��/�9O�]��� k����!������ s!�C�9�g�]�o�� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�??X� j�|ώϠϲ������� ��O�0�B�T�f�x� �ߜ߮���������_ �%_>�P��t��� �����������(� :�L�^�p�����c�� ������ $6H Zl~����� ��� 2DVh z������� 
//ן9�O/]����/ ���/�/ɟ۟�/?�� ??'?9?W?]?{?�� �/�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_?�X_ j_|_�_�_�_�_�_�_ �_�S_0oBoTofoxo �o�o�o�o�o�o�o� �,7�P�t�� �������(� :�L�^�p�����c�� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ����� �2�D�V�h� z�������¯ԯ��� 
���/9/K/a�o/�� �/}����/3��/ω? �?�?3�9�K�y�oϝ�����$MRR_G�RP 1���������  �`� � ������ @D7�  ��?������?������@T;g��Ũ���*�;�	l��	 �����X��'���F�O�^ �,X �k��Q�K��K���eK���K~o��K{GK�AM�sA�S��߈���?�;g?����@
���Р�����Iۿ�
���}v������X���4 � �p  �
�=ô7���A�� � >�L���=�������������Ѡ���(Ѵ��,  p_�  �����������������	�'� � )��I� �  {����:�ÈM�?È=���e���@u�{�v��������������ЈѸ����@�?��@�t�@���@�)��C6�B�O  CfK B�B���Q�����C�R�԰ � �_�� �ވ� H�B<�� ��a ����Dz��O��$J!�?�� �xy�jnz  ȅ:y��� ?�ff�ؿ��O ���,��8��/(*	�H��=$0(��V%P_(�z��U�UԿ�>�3�3����;��;�aʤ;r�@;���;�	�<�$D���/�A���+���?��� ?7fff�!?&02�A�5@�,%5iq1�-�� ]?��|?�'A���?�? �?�?�?�?OOAOSO0>OwOhF5F� fO �ObO�ON?�Or9�O+_~�HD�� E�J ���E9� E�0 4_m__j_�_�_�_�_ �_�_o�_oEo0e���nm2o�o�O�oXH)��C`5����t�Ɖ� EO�+8Ƈ�B�'o $6�*:��G?���_s9�B��@������yA� A��t<�	���@�7��[�F����d��k�����1��<��k���C����` Ca���j~��~�}�!�� �5��CH�f�CW�FB��1B-v�=����%������XR���u����z����ę�����AP���Blz��X���}�sp��R�d��
Ák�BU(�������F<rѵ���JGp@K���H�� I%�K�Ab!��L)-�yL!�GKӕ�#HP� H�R�����(�L&���J�3$H����H���A� �|�j�U���y����� ֯�������0��T� ?�x�c�������ҿ�� �����>�)�b�M� _Ϙσϼϧ������ ���:�%�^�I߂�m� �ߑ��ߵ��� ���$� �H�3�l�W�|��� ����������2��`/�h�S���w�G�E*<��~�C�?ټ����Ć�����CV���L7��\]G���_�(�Ya�`��,�%��<��1V��A3>�!3A��vM_�ܟv3�g�y�!��;�%D93�������	/��-/,�C P�"P_.na{o�/��/�/�/�/�+��/�/(?D?8<�8?G?V 8"�ta?#?�?�?�?�?�?��/mo'OOKO9K�`QO[O�OO�KO��O��O  �e 3��O�O__9_'_]_�kZ  2 D�f�EVp�U�Z�1B
��q
�C��Aj@��_jϜ�_~lD� D�ϕ�_>n|S�_�_zo�o�o�oj?� �aZ��UTjjXQrjyVZ�
 �o ,>Pbt�� ������[��a� ��I̿���Ld��2A� �@D<�U�?%`]� �� `��a�jA�XU�Ij��;�	9la�\!������xe�VPF��������5��'�VP#C� �P�����_� �?����ǟ���P���`��V_�z&'��9�pG���k���+UUp�s�=��ͭ���	�`Ϡ,bۯ�
�&f����G�TY3�֞u0 C '  [�e�:��-o A�[���u%b��ҿb��B�P�� @�Q.�abCp!��Tϛ� x�cϜχυ�j��.��  �j:v�a�`x#a���
�߮� R�d�
��0yߋ�>Ρ+`��
�����쿢>Lס �
��A����4��e%a�G�a�*�?fff?-�?&g��σ�&ib� �
�]���[���L桄 x����5� �Y�D�}��h����������_ F�P����7��X ��*�&���� ���-Q<u `������N /r;/�_/q/�/�/ 4�/�/V/�/�/?�/7?"?�R�_4�Qn� ,?�?|=(�0�~?�?�? O�? O9O$O]OHO�O lO�O�O�O�O�O�O�O #__G_2_k_V_h_�_ �_�_�_�_�_o�_1o Co.ogoRo�ovo�o�o �o�o�o	�o-Q <u`����� ����;�&�8�q� \���������ݏȏ� ���7�"�[�F��j� ������ٟğ���!� �E�0�i�{�f����� ï���ү����A� ,�e�P���t�����ѿ@�ο��+�R7(�����M�_�I�� mϣϑ��ϵ������� !��E�3�i�Wߍ�{�J�5P%�P����4 ���B����	�B�-� f�Q��u������ �����,��P��߹ ��������������� ��B0Rxfp����  2K� �*<N`r���������/"/A�F/T*
 T/N7�ߓ/�/�/�/ �/�/�/?#?5?G?Y?�k?��t/��{J���4�� ���1 �@D�  �1?�>�3 � `?7 �27 A�X�5���?� ;�	l�2��}��KC�0"K� F�����?/.�?:&�uO�L� �8�ObO@/ �O�O_�O%_]�0@�J_XW�x_��A���_�X_�_U+UU<�_�_=���ok�iS/`�09oGhjR&f�]oom�2�	�o6^u0  '�o�h�_�o�_x,�2ZO2�hBy Px~ @�`�u�aEC���o��o �����R�p&�.4�  ��r:h&Nq	~U�2�|j�|��� �в�ċjQ8�pڏ�>.a�0�1�z02�$�L�">L7a�jPA�=���;����s��2�3�2�p?fff?�p?&ǐ�� �t�2�4�y�5��8 =���D؟q�\����� ����ݯȯ����7���Ffp&�s�"� �����2���뿆�� ��3��W�B�Tύ�x� �Ϝ���������~_,� ��S߮�t�ҿ��߿� �����ߔ�
���O�`:�s�^���AfpA��������� �ꈕ�o��?�*�c�N� `������������� ��);&_J�n ������% I4mX��� ����/�3// 0/i/T/�/x/�/�/�/ �/�/?�//??S?>? w?b?�?�?�?�?�?�? �?OO=O(OaOsO^O �O�O�O�O�O�O_�O  _9_$_]_H_�_l_�_ �_�_�_�_�_�_#oo Go2okoVoho�o�o�o �o�o�o�o1C.�gR�vw(������{���� �'��7�9�K���o������ɏ���ی�P��P�Y��~O� �xT�~�i�����Ɵ�� �՟����D�/�h� S���w���W���=� �� �6�$�Z�H�~� l�������ؿƿ��� �.�  2��T�f� xϊϜϮ����������C�(�:�L�^�p�p�ߡ��ߴ�
 �� ��������)�;�M� _�q�������������{J������� @D��  �?�� �� `?��!��A��X��I� ;��	l!��}��k�e�%����F��a�K��������� ���=�����=( aL�p�y��0�������8z+v+UU03=���m��0���&f�������u0  '/'(K/vo/`��.���/Z(B �/�. @[ �%[!EC0�_/?[/8?#?�\?G?EO0�?�7 K �O2:�֮!
��!�W<�?�?n? !�O$K�8O0:OHJ>��)�M:�?�O��/��>L��� A���O�?�O�?O3!���!�� ?fff?� ?&'PR?C_O4.� "Q.�M9�}_��_V a�8_�_�_�_�_oo =o(oaoso^o�oR]`F� �o�o�o�on_ �Y�oK�ooZ� ~������� 5� �Y�D����R��� ԏ2��n��1�C� U��Oj�|������ӟؾ����A� A���'�0��T�?��E �>�����ï������ ���A�,�e�P��� ���������ο�� +��(�a�Lυ�pϩ� ���ϸ������'�� K�6�o�Zߓ�~ߐ��� ���������5� �Y� k�V��z������� ������1��U�@�y� d��������������� ?*cN`� ������) ;&_J�n�� ���/�%//I/ 4/m/X/�/�/�/�/�/��/�'(y���� ?;	???-?c?Q?�? u?�?�?�?�?�?O�?�)OOMO;Lv�P�BPN��{��/�O8�O �O�O_�O&__J_5_ n_Y_k_�_�_�_�_�_ �_o�Oy�Co��LoNo `o�o�o�o�o�o�o �o8&\J�jw  2o������� �2�D�V�d� ���������Џ�o��
 ��]O S�e�w���������џ������+�{B4����{J��$MS�KCFMAP  �-�� iwvD�E�  ]��ONREL  �qEt�jp]�EX_CFENB��
r������FNCƯ��JOGOVLIM���d����d]�KEYꦧ��_PA�N��-�)�]�RUN���]�SFSPDTY�@Ȧ�����SIGN����T1�MOT���]�_�CE_GRP 1-�-�t�\��	� �-�?ϗOc��sϙ� PϽ�t϶��Ϫ��)� �M��q߃�jߧ�^� ����������7��� [��P��H��l�]�QZ_EDIT���n���TCOM_C_FG 1�j����)�;�
��_AR�C_âqE�UA�P_CPL_�դN�OCHECK ?=j� pE�� ���������� 2 DVhz�������NO_WAIT�_L����װNUM_RSPACEg��wr=�7A�$OD�RDSP^�ѨO�FFSET_CAqR����tDIS��rPEN_FIL�E���=���SPT?ION_IO#�5���M_PRG %#%$*/".�WORK �緍ԣ G@S%��:mDC� ��m 9��m!	 ���m!�<����TRG_DSBL  -�Ᵽz��/��ORI_ENTTO����C���s�A rUT_SIM_D��q�D�TVXLCT �#B�@-5�_PEXE�g6RATs0	�ѥx�k2y�UP �<>%��.���?�?�?OI�$PARAM2�����}�&3	 d�� VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_���_ �_o#o5oGoYoko}o�o��<�_�o�o�o�o &8J\n��}�x����� � ��  ��  A�  B�p���B��3�pH>�p�  ���p�p+B�pp�p� 0�!�(�P Dz  �E;� E@ 7D���C� 0� �q����p�������)�+���r �E/!�,��qc�p���@�����_���#E	��C�/���/���������q���EZ�n�H� ���uL��� E�qX�J�L��t���;�D�p� ���`n�L�c�p���� ғ ����p�d������ d�� �(�:�L�L��qE� ��������  ���ҧL�Я��q� �(�:�L�^�p�����L���� �o���p��3���!�πD�R�ĽĽ���p� � '�Ϧϸ������� �.�DO]�o߁ߓߥ� �����������#�5� G�Y�k�}������ �_������1�C�U� g�y������o������ ��	-?Qcu ���#1�x��0� �}�<�*<N `r������ �//&/�J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?9/�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O i�˿ݿ�O�_%�_ M_[��OϘ_�9�� �_�_�_oo/oE�^o po�o�o�o�o�o�o�o  $6HZl~ ���������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v�������� �����?�*�<�N� `�r���������̯ޯ ���&�8��\�n� ��������ȿڿ��� �"�4�F�X�j�|�K� �ϲ����������� 0�B�T�f�xߊߜ߮� ���O�O��_C_)�7_ 1�[_m_�ߘ���-o�� ����������Eo�� p���������������  $6HZl~ �������  2DVhz�� ������
//./ @/R/d/v/�/�/���� �/۟�/��?*?<?N? `?r?�?�?�?�?�?�? �?OO&O8O?\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_KO �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o{����C�)7� !_m��o��-�?� )������A��q��$PARAM_�GROUP 1��gX��oL�`8� � ��q��� @D� M ��?�����?�p����qC>�����t~�  ;�	l���	 �����X��΀π���^ �?,X ���p�H��H�ff�H�  H���H�WH-����|�#�o�oi���qB��  B��������������s�4  ��p  �
=É��������ȟ��sA�8�¼r=��q«�C���r,�2���G��wρ[���|,  � _�  ������M  Д������u	'� � �ТI� � � ��l�=��q������@�@"����F�������[�i�2���������-CݐB���f�������б��Ŀֿ�   ���CR>���� :��<�H��wB�L�+�Xŷ�c 3�tŕqDz�������Ϧ�����Ȯ?�� �x ��n!�  �,�:˅��!D� ?�f�f{R�d��� ���ߪ���8�����ڐ��D�����(����P��!�A�����f�>��33}���;���;aʤ;r�@�;��;�	��<$D4�q��A)�s봂��?3�q�o?fff��?&�����A���@�,����©ᵄ�� �����#���脃�X� C�|�g����������� ����0T?x�����q�mD��� E��j E9� E�0�& J5nY�}� ����{�-�:/ �[/��/��/�/�/x�/{���?��|�3��BA��/=?(?a?hL?�?p9A+�A�4 㠰1�?��y?�?u?O�<?��OOKO�6OaI���k^OC}����` Ca[O�H*%D�%@$A�A@I��ܾ��CH�f�CW�FB��1B-v�=����̞������XR���u��!_DA�ę�����AP���Blz��X���$_0��R�d��
Ák�BU(�������E@K����JGp@K�ÌH�� I�%K�A	�aLL)�-yL!�GK���#HP� H��R��_�P(�L�&��J�3$H�㞀H���A��_#_o�_5o oYo Do}oho�o�o�o�o�o �o�o
C.Sy d������	� ��?�*�c�N���r� �������̏���)� �M�8�q�\�n����� ˟���ڟ���#�I� 4�m�X���|�����ٯ�į֯���3��G�x��b�%�C�?�c��j�Ć�����C�V�������޿����O�:�s�^Ɲ(d��`���0��y���dų1V��<��^�3>��������v��߰?�v3�g� �2��!�;�%D93ҵ�L�Lٌ�z߰�p������^� Pl�	P�!"//��;�0e�P��t���������������8�0t���S�>�w�b����B�/������������8&HO��HZ  �e 3�t6�����  2 D��7E� 1�b��B�1�1�0C��@
��A��@�?z��~�D� D��������/!/3/�E/W/��?�p!��J������oA��9 ��
 ^/�/ �/�/�/	??-???Q?�c?u?�?�?�?���! {����̿���ӀK�&��1 @�D�0�1?vPA � `V�By��4�1��2L;�	lBᖃ�RKLC@iK��F����2O�?�O��1��O�L��C��O�O���i&_��J_5_n_ Y[]`@�_�W��_!��A��_�Xa_o]U�+UUoo=���Tofk cv`�0�o�hb&f�o�m�2�	�o>}^u0  '��v�A�D,W_Pb K�B�OyAxBU��| @e�t4C�F�B�
�C��.�,b6�m�{�  �6�:�"�!� ��B>���ÏU� �����=�+� �2�>ua�0V�=�y�k��FI�>L~a�T=�A� ����ۏi%	A�3B��p?fff?�p?&�9�*�6�B	�&} �Ed�H���HD� ����ܯǯ ��$�� H�Z�E�~���g����� ؿO�q�s�ѿ2�ͿV� A�z�eϞωϛ��Ͽ� ������@�+��_s� 9ߚ��������U�� �*�<�۟Q�c��ߖ�������T� �Q_��8�#�ϕ�o %���q����������� ��(L7p� m������ �H3lW�{ �����/�2/ /V/A/z/e/w/�/�/ �/�/�/�/??@?R? =?v?a?�?�?�?�?�? �?�?OO<O'O`OKO �OoO�O�O�O�O�O_ �O&__J_5_G_�_k_ �_�_�_�_�_�_o"o oFo1ojoUo�oyo�o �o�o�o�o�o0 T?x�u���z�w(�q���� ��&��J�8�n�\� ~�����ȏ���ڏ�P��4�"�]�P̒Pf���b�����x��ş ���ԟ���1��U� @�R���v�����ӯ�� ����`�*���3�5�G� }�k�����ſ���׿�����C�1�g�u�  2�ϭϿ�����@����+�=�K��� o߁ߓߥ߷��������
 ����D�:� L�^�p������������ ��b����7{J�_�+�[��H� @D�  �\�?�b� � `?��h���C]�\�X�>�� ;�	lh�c�}�����l�����F�������+����.�Є�N	 �߄o����]������]�Y�.��@N�r�+UyUwz=��ʹ��`�X���a&�f/-N�[�:/�u0  '`/n(a �/��/�u��/�(�B �/> @� 45�!ECw��/[?@�/?j?�?�?��0\�?�7  Ȗ2:�$S��!%h��<O#O�? .�YOkK"�18�0�O�J>�I��p�:�?�O�/)�>L�Sĝ0A��ODO�O�<O�3h�N�h�10?offf?40?&nP �?�_�4u�iQu��9d� �_b��_SV��_oo <o'o`oKo�ooo�o�o �o�o�o�o�o8�_ �_�_1�-��� ����4��X�C� |�g�����%ӏ���� U�yB���f�x��� ��;_��ß]�������>�)�A0A�f��n�w�6�����/U 7/���ѯ
����@� +�d�O���s�����п �Ϳ��*��N�9� r�]�oϨϓ��Ϸ��� �����8�J�5�n�Y� ��}߶ߡ�������� ��4��X�C�|�g�� ������������	� B�-�?�x�c������� ������>) bM�q���� ��(L7p �m������ /�/H/3/l/W/�/ {/�/�/�/�/�/?�/�2?7($1��� T?f;P?�?t?�?�?�? �?�?�?�?(OOLO:O�pO^O�O�L��P,RP�N Q¤%?�OI8�O %__I_4_m_X_�_|_ �_�_�_�_�_o�_3o oWo�O���o䈓o�o �o�o�o�o%I 7Ym����w  2Ro���1��C�U�g�y������� �Ϗ����)�HoM�[�
 [�9��O ������П������*�<�N�`�r��B{��o�{J��������B�� @D� � ��?�£ � #`?>�Ȣ>�C����|�F� ;�	lȢ�A}���̠)�E�F����6���A��|���E�䨮� i�G��Ͽ��,�� �� �Q�_ǽϹv���РϮ�!����+�UU����=��� �&���6и�@�N���&fd�vݮ��y��=�?u0  '���� �������բa�9���B W�� 1@����EC�A��������������-�;�  ���:Ho��qU��uȢ��8q���� �@��D����8������>5р��С��9�+S>1L>ѳt��A�D��B����Ȣ��Ȣ���?fff?��?& � �����բ�դ�� ĥ$¨D���x c������/ //>/P/'/t/_/�/ 13�/�/�/?? :?%?^?I?[?�??�? �?�?�? O�?��3O�? ZO�/{O�/�OO�O�O �O�O�_#_�OV_A_�z_e_�_�_Am�A��T��S�_�_�_�Z ����_Fo1ojoUogo �o�o�o�o�o�o�o 0B-fQ�u� ������,�� P�;�t�_�������Ώ ���ݏ��:�%�7� p�[��������ܟǟ  ����6�!�Z�E�~� i�������دï���  ��D�/�h�z�e��� ��¿���ѿ
���� @�+�d�Oψ�sϬϗ� ���������*��N� 9�r�]�oߨߓ��߷� �������8�J�5�n��Y��}�(��������������
��� .��>�@�R���v���@����������eP�	P&=A"d��V�� [�p����� � K6oZ �~�^ O�DH� �/=/+/a/O/�/s/ �/�/�/�/�/?�/'?7  2�[?m?? �?�?�?�?�?�?�?JJ?/OAOSOeOwO�O8��O�J
 �O�G �O__0_B_T_f_ x_�_�_�_�_�_"�O���{J��$P�ARAM_MEN�U ?�U��  �DEFPULSE��[	WAITT�MOUT/kRC�VBo SHE�LL_WRK.$�CUR_STYL�-`nlOPTAL9a�oTB�o�bCioR_DECSN:` �l�o�o1,> Pyt�������	�aSSREL?_ID  �E1���USE_PR_OG %j%�j��CCRF`*�1�c}�_HOST !j!����w�AT7 ��ۃ����݃|�v�_TIMEDb�*���`GDEB�UG(�k�GINP_FLMSK@��o�TR~� q�P�GA�� _��I� ���CH}�  �q�TYPEl@��4�]�X�j� |�������į���� �5�0�B�T�}�x��� ��ſ��ҿ���� ,�U�P�b�tϝϘϪ������q�WORD �?		FO�LG-c	U�	�MAKRO+�S�UCHL�C2�S�7T�TRACEC�TL 1��U�a
 0[ \~�@ � �{��2�ߗߩ�S�DT� Q��U��o��D �  U��������T*���������U��������U��������T�@��������Tސ��!��"��#��U$��%��&��'��U(��)��*��+��U,��-��.��/��U0��1��2��3��U4��5��6��7��U8��9��:��;��U<��=��>��?��@�Ԙ`�Ұ`���`��'���-`��F��\���H��I��J�����B���M���`��6���D7 ��Q�ԝ���S��TF`��U��V��W��UX��Y��Z��[��U\��]��^��_��U`��a��b��c���d��e��f��	��ϐ ) ®��) ��ĳN�r���1��P���z������T��	�
��	������ "� �*� 2g h�On�g j�����	Pql�Qqn�co�R�Sqq
�T�T������g s{́bR�U��U�U�@��
�f�ԭf��	_�_�_*�_$_)$_G ��G R_Y_1f�	�f�f�f!�	U`�`�`�$��$�$�&�$$�	$$�$!$�)$1$9$��$�I`$`!$`	fV1�	a�a�a��a$a!$a	1� �s�s�sJ�����6������6�	�!J)19��)�U)�)�)�)��)�� g��������������������������������������������������������������������������������������������
 .@Rd�o�]C�is��g�m��� //$/���ԆA$���d��d)$�q$y$�$Y�d�	���*!�f�Tf�Tf�/�/��/�/?#?577 �Sf��Tf�T�Y4���d��d�d6�;����;q����e��2�r��)��)���)��)��)��)��)	�)�)�)�!�))�)1�)9�)�A�)I�)Q�)Y�)�a�)i�)q�)y�)���)��)��)��)���)��)��)��)���)��)��)��)���)��))	)�))!)))�1)9)A)I)�Q)Y)a)i)
q)y)�'A�5o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{��5 k�����% 7I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_o#o5o GoYoko}o�o�o�o�o �o��o1CU gy������ �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q����� ����˟ݟ���%� 7�I�[�m�������� ǯٯ����!�3�E� W�i�{�������ÿտ �����/�A�S�e� wωϛϭϿ������� ���o=�O�a�s߅� �ߩ߻��������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ������1CU gy������ �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?1�?�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y�����s?��ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� �������������� '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o��1o Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u���$PGTRACELEN  v��  ���A`ȋ�_UP ������������y����_CFoG �����*Aa������ĝ�����������DEFSPD ����@a��Ћ�IN~��TRL ������8��V�PE_C�ONFI�����O�����#�WLID�á���ԿGRP 1���� �v�CH�����Aa�A�  G�G �G�7�F�, A�  D	���A`d��)�9��?� 	 ����S� ´��n��B���������������B>��e�G�Y�C� <,?1<49X^��� Z�����������v� @9��IoZ�z�����
 C��f��.X��A�NB�RH[���HL�rG/"�����=�(Ms^  >W?�>V��z�@v���/^�!���
V7.10be�ta1� @��33@2�\@�;�CRA`C C_>  CW��T#/D�� j"0�g!~�D�� Dj\ �2 ��B�\ S C�] �p���!~���CRp�B���B ��@��� h� A �]�� `ffA�����T"���/?����&�8�ѩ� �[?�?j?�?�?�? �?�?�?�?!OOEO0O iOTOyO�O�O�O�O�O �O_�O/__,_e_P_ �_ܳ �_�_n_�_�_ �_oo=o(oaoLo�o po�o�o�o�o�o�<./T#F@ >y:}N`|~ ?�&� �����/�??/? A?J��on���k����� ȏ���׏����F� 1�j�U���y�����֟ �ӟ���0��T�?� x����_����o��ϯ ��,��)�b�M��� q�����ο���� 1c=�O�y���� �������	��-�?� H��l�Wߐ�{ߍ��� ���������2��V� h�S��w������ ������.��R�=�v� ������[������� ��*N9r�o ������/� a�;Mn�ϒ������$PLID_�KNOW_M  }:%�>!~�SV ���v������)/;/M/�q/\/�n/�/�� �M_?GRP 1��� �lCR�"��� �&�$ �z0H��@�( "1*5&?8<���	7�+ a????�?S?e?�?�? �?	O�?�?9O�?OuO�+D�MR�#��-T���C5��"�C� � ��O�N_�O�� �O>___$_�_H_�_`�_~_�_�_�%ST�!�1 1��"`�> 0EZ!�D��f��.X���ANB�RH�[��HL�rG�/"����Fvo  [omoo�o�o�o�o �o�o!bEW��{����m2o)`� �C��8� J�x�n�����ӏ��ȏ ڏ����"�c�F�X��j����������k3 �(��̟-�n�Q�c� �������������� 4��)�;�M���q��� Ŀ������c4�'� �˿,�m�P�bϣφ� �Ϫϼ�������3�� (�:�Lߍ�p߂��ߦ�(����c5�&��'�<)�n6�%�7�I�c7b�t���c8��������cM_AD  �$"c�  dPARN_UM  ��"��!��7�T_SCH
N� \�
��o�����UPDo����?S_CMP_� Q����'�S_E�R_CHK6����cO3ERS8�@��"_MOP���_��RES_�G`�� ?aDA��lB�&I�,c�G@F �OOUL16gZ� ~�����	/� -/���1//�/y/ �/�/�/�/�/?�/(? ?L???Q?p?6/�� Q/�?u?�?�?	O�?-O  O2OcOVO�OzO�O�O �O�O�?���?�O�O D_7_h_[_�__�_�_ �_�_�_
o�_o.o�O��\_Qo�a� no�o�o���o�o�o�����o�V �1����� ��^�`�^h�]�T�]���THR_INR� �S��d�d�vMA�SS� Z�wMN���sMON_QU?EUE �š���ȡ�%MJ� �2��y��4A��  @�߉�Bʪ��!	�N- U�qN�v_m�END8o����EXE�������BE��y�j�OP�TIOv��m�PR�OGRAM %��z%l�J3�k�T�ASK_IP�ߎO?CFG ��|����ODATA��1�}�@  ��) 2 gޟ���&�0��ڑ i   �, 6 ? G R ^ gF�X�j�H|���C�"����௯��ӯ��� ����ڟ*�<�N�`�4� ����������̸C����� ��$�6� ����j�|ώϠ�t� ȿƿ��������5� 1�C�U�g��Sϣߵ� �����߿���!�3� E�+�y�{����s��INFO���}���#
��.�@� R�d�v����������� ����*<N`�r��I���� �=is���DIT ��}�@mU����WE�RFL��rs��RG�ADJ �}�A�  '?��3�q�m�x��U��?C�ѐ <@�����%qq����I�J��U˒5��\9fqrb�bA<t�t$&�* /" **A:""��/'#UL"FG%��!Q)Q� ��q/sE/W/i/{/�/ �/�/�/�//?�/?? �?�?S?e?w?�?�?�? �?�?�?�?OO+OUO OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ �_�_�_�_�_$o�_�_ �_oko5oGoYo�o�o �o�o�o �o�o�o ;1CUg��� �����	��-��?�Q�c�u������ 	��,��P�;�	)u� #A���=�Ɵ��� 
//�@/ʏ܏q� � ��L�^�˯�������� �ܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�Dϱ�h� zόϞ���������� N��.�@߭�d�v߈� ������������ *�<�N�`�r���� ����������&�8� J�\�n����������� ��G��"4�X j|����
C .l�v<�8�؟ ���� �2���� ��>/P/b/t/�/�/ �/�/�/;?�/??(? ~?L?^?p?�?�?�?�? �?7O�? OO$ONOHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_o�_�_�_ 
owo.o@oRodo�o�o �o�o�o�o�os *<N`���� ������&�8� J�\�n��������#� �G�^h����R��� ş�� /*/�6/�� ҏg�����B�T�~�x� ��������ү���� �,�>�P�b�t����� ����ο�M���(� :ϧ�^�pςϔ��ϸ� ����I� ��$�6ߣ� Z�l�~ߐߺߴ����� ����� �2�D�V�h� z������������ 
����@�R�d�v��� ��������&�� �<N`r����  9Kb�l����.���$PRG�NS_PREF ����� � 
�IOR�ITY  ݔ�����MP�DSPON  `ݖ���#UT&��5&ODUCT_�ID �"���OGGRP_�TGL$m&V&TO?ENT 1�i*��(!AF_IN�EE �/�!t�cp�/�!u�d�/�!ic�m!?�Z"XY_�CFG ��+ ;��)� #��?�?� ��?�?�5�? �?�?!OOOWO>O{O bO�O�O�O�O�O�O_i*Y#t3�� %�xO_a_�?#O~��#�/�:_�_���-%�X�A���,  ���_
oo.o)(T����0"��PORT_NUUM#� %��_CARTREP�& {<�SKSTA�E' �jSAVE� �i*	26�00H601��!�_'3?KC 	ox����ݓe������
��|JU��e_�  �1��+ p �4R����#��������a_CONFIw0�Zg#�]�U��ޔ��0����ȃPt22�֋���[���C�U��$�q�2��։�a����Z8��T�����+���C���:?~��^�k�?���ۏ��U��Dt�,?1DL������ɟ)#ݑ?�k\���p�� �� ��ݑ�y���i��� ��_������_��U]� �A���Q�w��ۯ�� ���#����Y��=� ˿)�sυ�׿鿻��� ����U���9�Kߝ� �ρߓ��Ϸ������ ����c߭�G�Y��}� ���ߛ����)�s�� ���C�U���y�����~k2S_MOTI$ ;2�֋
�?����_��);M��`�5����x�<l�Z+= Oas����� ��y��#�&/./ @/R/d/v/�/�/�/�/ �/�/�/:�/7?I? [?m??�?�?�?�?�? �?�?O
??EOWOiO {O�O�O�O�O�O�O�O __/_*O<Oe_w_�_ �_�_�_�_�_�_oo +o=o8_J_Jo�o�o�o �o�o�o�o'9 K]Xojo���� ����#�5�G�Y� k�fx���ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����������)� ;�M�_�q��������� ��Ư���%�7�I� [�m�ϑϣϵ����� Կ��!�3�E�W�i� {ߍߟ߱��������� ���/�A�S�e�w�� ������������ �=�O�a�s������� ���������"� "]o����� ���#50B k}������ �//1/C/>Pb �/�/�/�/�/�/�/	? ?-???Q?c?^/p/�? �?�?�?�?�?OO)O ;OMO_OqOl?~?�?�O �O�O�O__%_7_I_ [_m__�_�O�O�_�_ �_�_o!o3oEoWoio {o�o�o�o�Q�Q�Q�e��i%�f�o�fEL <�o  '��m�c<�S�e  8R�Q8_���� �_�_� 	��-�?�Q�c�u��� ������Ϗ�_��� )�;�M�_�q������� ��˟ݟ����%�7� I�[�m��������ǯ ٯ�����
�
�E�W� i�{�������ÿտ� �����*�S�e�w� �ϛϭϿ�������� �+�&�8�J�s߅ߗ� �߻���������'� 9�K�F�X߁���� ���������#�5�G� Y�T�f�x�������� ����1CUg yt�������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ ���/�/??%?7? I?[?m??�?�?�?�? �/�/�?O!O3OEOWO iO{O�O�O�O�O�O�? �?�O_/_A_S_e_w_ �_�_�_�_�_�_�_�O _+o=oOoaoso�o�o �o�o�o�o�o�_o "oK]o���� �����#�0 Y�k�}�������ŏ׏ �����1�,�>�P� y���������ӟ��� 	��-�?�Q�L�^��� ������ϯ���� )�;�M�_�q�l�~��� ��˿ݿ���%�7� I�[�m��z������� �������!�3�E�W� i�{ߍߟߪì����Ղ��%��������� ��%���Ӡ��� � (�B��8�O����� �Ϯ������� /�A�S�e�w������� ��������+= Oas����� �����'9K] o������� ���5/G/Y/k/}/ �/�/�/�/�/�/�/? //C?U?g?y?�?�? �?�?�?�?�?	OO? (?:?cOuO�O�O�O�O �O�O�O__)_;_6O HOq_�_�_�_�_�_�_ �_oo%o7oIoD_V_ h_�o�o�o�o�o�o�o !3EWidovo �������� /�A�S�e�w����� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o�����������ğ� ���#�5�G�Y�k�}� ������ſ��үҿ� �1�C�U�g�yϋϝ� �����������-� ?�Q�c�u߇ߙ߽߫� �������� ��;�M� _�q��������� ����� �I�[�m� ��������������� !�.�@�i{� ������ /A<Nw��� ����//+/=/ O/a/\n�/�/�/�/ �/�/??'?9?K?]? o?j/|/�?�?�?�?�? �?O#O5OGOYOkO}O@�O�3�1�1�E�I%�F�O�F���O�O�Ox�E�3�E  _2_�18?_u_�_>�_� �?�? �_�_�_oo1oCoUo goyo�o�o�o�?�_�o �o	-?Qcu ������o�o� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ�����
�3�E� W�i�{�������ïկ ������*�S�e� w���������ѿ��� ��+�&�8�a�sυ� �ϩϻ��������� '�9�4�F�Xρߓߥ� �����������#�5� G�Y�T�fߏ����� ��������1�C�U� g�y�t��������� ��	-?Qcu ��������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ ���/�/?!?3?E? W?i?{?�?�?�?�?�? �/�/OO/OAOSOeO wO�O�O�O�O�O�O�? �?O+_=_O_a_s_�_ �_�_�_�_�_�_o�O _9oKo]ooo�o�o�o �o�o�o�o�ooo 0oYk}���� �����1�,> g�y���������ӏ� ��	��-�?�Q�L�^� ��������ϟ��� �)�;�M�_�Z�l��� ����˯ݯ���%� 7�I�[�m������������%����ʹ��� ~h���������  �"ς�8�/�e�wω�� |��������� ���!�3�E�W�i�{� �ߟ�r���������� �/�A�S�e�w��� ����������+� =�O�a�s��������� ��������'9K ]o������ �����#5GYk }������� �C/U/g/y/�/ �/�/�/�/�/�/	?? /(/Q?c?u?�?�?�? �?�?�?�?OO)O$? 6?H?qO�O�O�O�O�O �O�O__%_7_I_DO VO_�_�_�_�_�_�_ �_o!o3oEoWoiod_ v_�o�o�o�o�o�o /ASewro�o �������+� =�O�a�s������� ͏ߏ���'�9�K� ]�o������������� ����#�5�G�Y�k� }�������ů��ҟ�� ��1�C�U�g�y��� ������ӿί��� -�?�Q�c�uχϙϫ� ��������� �)�;� M�_�q߃ߕߧ߹��� �������� �I�[� m����������� ���!��.�W�i�{� �������������� /A<�N�w�� �����+ =OJ\���� ���//'/9/K/�]/o/z|r�%�)%8�&�/�&�/�/�/�%p�%  8�/?r8?U?|g?y?� l ~�?�?�?�?�?O#O 5OGOYOkO}O�Ob�? �O�O�O�O__1_C_ U_g_y_�_�_�_�O�O �_�_	oo-o?oQoco uo�o�o�o�o�_�_�o );M_q� ������o�o� %�7�I�[�m������ ��Ǐُ���
�3� E�W�i�{�������ß ՟������A�S� e�w���������ѯ� �����&�8�a�s� ��������Ϳ߿�� �'�9�4�F�oρϓ� �Ϸ����������#� 5�G�Y�T�fϏߡ߳� ����������1�C� U�g�b�tߝ������ ����	��-�?�Q�c� u������������� );M_q� �������� %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ ���??/?A?S? e?w?�?�?�?�?�?�? �/�/O+O=OOOaOsO �O�O�O�O�O�O�O�? �?O9_K_]_o_�_�_ �_�_�_�_�_�_o_ _GoYoko}o�o�o�o �o�o�o�o1,o >ogy����� ��	��-�?�:L u���������Ϗ�� ��)�;�M�_�j�l��b�x���%s�����N� ]��͟ �{�����`���  8��b�8�E�|W�i�� \� n�����˯ݯ��� %�7�I�[�m��R��� ��ǿٿ����!�3� E�W�i�{ύϟϚ��� ��������/�A�S� e�w߉ߛ߭ߨϺϺ� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ��������������# 5GYk}��� ������1C Ugy����� ��	/(Q/c/ u/�/�/�/�/�/�/�/ ??)?$/6/_?q?�? �?�?�?�?�?�?OO %O7OIOD?V?O�O�O �O�O�O�O�O_!_3_ E_W_ROdO�_�_�_�_ �_�_�_oo/oAoSo eowor_�_�o�o�o�o �o+=Oas ��o�o����� �'�9�K�]�o����� ����ۏ����#� 5�G�Y�k�}������� ����ҏ����1�C� U�g�y���������ӯ Ο��	��-�?�Q�c� u���������Ͽ�ܯ � �)�;�M�_�qσ� �ϧϹ���������� �7�I�[�m�ߑߣ� �����������!�� .�W�i�{������ ��������/�*�<� e�w������������� ��+=OZ�\�R�ht	%c��y �� � �txtP�t  ��R�8�5G>Y� L�^� ������// '/9/K/]/o/B�|�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�/�/�? �?�?�?OO1OCOUO gOyO�O�O�?�?�O�O �O	__-_?_Q_c_u_ �_�_�_�_�O�O�_o o)o;oMo_oqo�o�o �o�o�o�_�_�_% 7I[m��� ����o�o!�3�E� W�i�{�������ÏՏ ������A�S�e� w���������џ��� ���&�O�a�s��� ������ͯ߯��� '�9�4�F�o������� ��ɿۿ����#�5� G�B�T�}Ϗϡϳ��� ��������1�C�U� g�b�tϝ߯������� ��	��-�?�Q�c�u� p߂߂��������� �)�;�M�_�q����� ���������% 7I[m���� ������!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�� �?+?=?O?a?s?�? �?�?�?�?�?�?�/�/ 'O9OKO]OoO�O�O�O �O�O�O�O�O_OO G_Y_k_}_�_�_�_�_ �_�_�_oo_,_Uo goyo�o�o�o�o�o�o �o	-?JcLaBa�Xudy%Sv}�v�y�t� �
�d}xds@cdu  ��Ba8�%�7�>I�� <oNo ��������Ϗ��� �)�;�M�_�2ol��� ����˟ݟ���%� 7�I�[�m��z����� ǯٯ����!�3�E� W�i�{���������տ �����/�A�S�e� wωϛϭϨ������� ��+�=�O�a�s߅� �ߩ߻߶������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ���������1CU gy������ �	?Qcu �������/ /)/$6_/q/�/�/ �/�/�/�/�/??%? 7?2/D/m??�?�?�? �?�?�?�?O!O3OEO WOR?d?�O�O�O�O�O �O�O__/_A_S_e_ `OrOr_�_�_�_�_�_ oo+o=oOoaoso�o �_�_�o�o�o�o '9K]o���o �o�o����#�5� G�Y�k�}�������� ������1�C�U� g�y�����������Ώ ��	��-�?�Q�c�u� ��������ϯ�ܟ� �)�;�M�_�q����� ����˿ݿ����� 7�I�[�m�ϑϣϵ� ���������
��E� W�i�{ߍߟ߱����� ������/�:�<�2��H�T�%C�m�w�ocykd�� me=T�xT�0�T�  ����2�8���'�>9�� ,�>� w��������������� +=O"�\�� ������ '9K]oj|� �����/#/5/ G/Y/k/}/x��/�/ �/�/�/??1?C?U? g?y?�?�?�/�/�?�? �?	OO-O?OQOcOuO �O�O�O�?�?�?�O_ _)_;_M___q_�_�_ �_�_�_�O�Ooo%o 7oIo[omoo�o�o�o �o�o�_�_�_!3E Wi{����� ���o/�A�S�e� w���������я��� ���&�O�a�s��� ������͟ߟ��� '�"�4�]�o������� ��ɯۯ����#�5� G�B�T�}�������ſ ׿�����1�C�U� P�b�bϝϯ������� ��	��-�?�Q�c�u� pςϫ߽�������� �)�;�M�_�q��~� �ߢ���������%� 7�I�[�m�������� ��������!3E Wi{������� ���/ASe w������� //+/=/O/a/s/�/ �/�/�/�/�/�/�� '?9?K?]?o?�?�?�? �?�?�?�?�?�/?5O GOYOkO}O�O�O�O�O��O�O�O__����$PURGE_E?NBL  ,A-A��-A4PW}F<PDO  DT4,BOQ TR_I]TgQ�KUTQRUP_�DELAY ��"A"AKU,B�R_HOOT %�UiR%+B��_�]�SNORMA�L�XKR�_!o�WSE�MI o&oeopQQS�KIP_GRP �1ĞUMQ x 	 ho�o�o �o�o�o�i�U'w GYk1�}�� �����1�C�U� �e���y�����ӏ�� ����-�?�Q��u� c���������͟����)�;��U�$RB�TIF^T�ZY�CV_TMOUT^V�U��Y�DCR�cƾ�i ��a=���,AEd[e�B9�*,AB��|�m����h{0@ u��ӷ��o���;��;�aʤ;r�@;���;�	�<$D�/@�j�{� {�����ſ׿ �����1�C�U�g� ����vϯϚϿ����� 	�L�-�?߂�c�u߇� �߽߫��������� )�;���_�J��n�� ����� ���V�7� I�[�m���������� ����������3W B{f������ *�/ASew������,kRD�IO_TYPE � �[��RE�FPOS1 1Ǟ�[
 xSoY) �}/��/�-L/^/�/ �/�/?�/A?�/e? ? b?�?6?�?Z?�?~?O O�?�? OaOLO�O O �ODO�OhO�O_�O'_ �OK_�Oo_�__._h_ �_�_�_�_o�_5o�_ 2okoo�o*o�oNo�o��o/%2 1�;+ J/�o�oL�opvo� /��������6��Z�l�-'3 1�
��V�ԏ���� ����@�ۏ=�v�����5���Y��p�0$4 1ʍ�����۟Y� D�}�����<�ů`�¯ �������C�ޯg���0$5 1���&� `�޿ɿ��&���J� �Gπ�Ϥ�?���c�x��z�0$6 1�;+������`��τ��3!7 1��.�@��z�������S8 1α�������x����/�SMASK 1�� H ������XNO���4��D�/!MOTE  ��M�_CFG ��[�D�."PL_RGANGW�+!_���OWER �;%���g�."SM_D�RYPRG %�;*%X� ��TAR�T ���
UME_PRO����j�,$_EXEC_E�NB  �c�G�SPDC � �<e��GTDB��
sRM��MT_���T��Y��OBOT�_ISOLC����x'NAME� ;*KJ�BVTU2111�60R01xB �V#_ORD_N_UM ?��
!_H6�8��895  ��+!���������|� ��/ PC_TIME�OUT�� x/ S7232t�1�;%�� LTEA�CH PENDA�N�p�G�I�n�W��Maint�enance C�onso�C�R,"�b/��	UnbenutztY*�/X/�/��/�/�/�/�b"NPqO �K����SCH_LF ����	�1T;MA�VAIL��5���c�SPACE1 {2��
 K?@HHG�v�F�������4L8�?� L;WOL?;O�O�O�O�O �G�?OO%O�OIOkO ]_~_A_�O�_�Y�#� �]�O__%_�_I_k_ ]o~oAo�_�o�o�o�O �_o!o�oEogoYz =�����o�o /�Suw9��� ����������+� ُO�q�c��������� ��ߏ���'�՟K� m�_���3�������˯ ����#�ѯG�i�[� |�?�������ǿ��� ��1�C�U�WϾ�;� �Ϯυ������	�� -���Q�s�e�7߉ߪ��ߓߥ��52�?�?�� �#���G�i�x��\� ����������*�<� N�`�r�t���X����� ������&�8�J��� n����T���� ��"4F�j� ~�R���� 0B�f�z/�/ ^/��/�/�///,/ >/�/b/�/v?�?Z?�? �?�?�???(?:?L? �?p?�?�?VO�O�O�O �O OO$O6OHO�OlO �O�_�O�_�_�_�_�O _ _2_D_�_h_�_|o �oPo�_�o�o�o
oo .o@o�odo�ox�\ ������3��
� .@�d����� y�ˏ�ӏ�5�G� Y�k�}�������u�ǟ 蟿����1�C�U�g� �������q�ï��� ͯ�-�?�Q�c���� ������o����ٿ� )�;�M�_�σ����� ��{�ݿ�����%�7� I�[�	�ϡϓߴ�w� ��������!�3�E�W� i��߯߱�s����� �����/�A�S�e�� �������������� �+�=�O�a����� ��m����' 9K]����@y���/�4� '�9K]/���/ �/�/�/	?�/?#R/ d/v/�/�/�/�??�? �?O�?O<?N?`?r? �?2O�?�?�O�O�O_ _�O8OJO\OnO�O._ �O�O�__�_�_o�_ $oF_X_j_|_*o�_�_ �o�o�o�_�o Bo Tofoxo&�o�o�� �����>Pb t�4������� �ڏ�:�L�^�p��� 0���ȏ���ޟ��� ��6�H�Z�l�~�,��� ğ��ׯ�������"� D�V�h�z�(��������ӿ���	���#+52.D/V�h�z�(Ϟ� �����ϳ��&��;�#+6O�a�sυϗ�E� ���������"�C�*�X�#+7l�~ߐߢߴ� b�����	�*���?�`�G�u�#+8����� ������&G
\�}d�#+G �N5+ �:
�  �,: 5%K]o������ ��o�>d � %/7/I/<j/|/�/�/ ����*�/�+?
/ ;?M?_?q?d/�?�?�? �/�/�/�/?O7O*? [OmOO�O�?�O�O�O��?�?�?O$O6_ `� @> oU� }_�O�_�Ek_9_�_-O o�_�_�_�_loo1o So�ogo�A�a�E�c�o �o!�e�oSe �9k���������L
�_n�@��_MODE  ����S ��]�_Z���_��9�	4�]�D�CWO�RK_AD���{��F�R  ����b���_INOTVAL��������R_OPTION�̖ ��F�TC�F� ۗ���?���7���V_DATA_GRP 2��H�DU@PJ�y�F� ����G�ʯ���ܯ�  �6�$�F�H�Z���~� ����ؿƿ����2�  �V�D�z�hϞόϮ� ���������
�@�.� d�R�tߚ߈߾߬��� �������*�`�N� ��r��������� ��&��J�8�n�\�~� �������������� 4"DjX��Be� �������q�5 #YG}k��� ����//C/1/ O/U/g/�/�/�/�/�/ �/	?�/??-?c?Q? �?u?�?�?�?�?�?O �?)OOMO;OqO_O�O �O�O�O�O�O�O__ _%_7_m_[_�__�_ �_�_�_�_�_�_3o!o WoEo{oio�o�o�o�o ��o� ��o�oA we������ ���=�+�a�O��� s�������ߏ͏�� '��3�9�K���o��� ��ɟ���۟����� G�5�k�Y���}����� ���ׯ���1��U� C�e�g�y�����ӿ�� ����	��Q�?�u� cϙχϽϫ������� ��o>�b�M�ߕ� ߹ߧ��������� �%�[�I��m��� ���������!��E� 3�i�W�y�{������� ������/e S�w����� ��+O=sa ������/ /9/'/I/K/]/�/�/ �/�/�/�/�/�/�/5?�#?Y?+��$SAF�_DO_PULS�  -��������1t0CA?N_TIME�0}���3���1R ������8�		����
�8����4�4��  ^�OO0OBOTOfO�?��O�O�O�O�O�O�G��1  B2�T�1�1dXQ Q��4}��1�� @ CVT[�0P_z_�\�1�_��WP�U�� {@B�3T i_��_�_oiT D��oAoSoeowo�o �o�o�o�o�o�o�+=OaX^?VNV{py 
�q�p��y�3�1;��o}��4p{}
�t� �Di�0��A�1�z�� ��B�1�q�1�A�1�z�Y�k�}�������  ��������  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v���������@Я�����$��h_ H�Z�l�~�������ƿؿ'�>T�Q���R �7�I�[�m�ϑϣ�Žρ�0�22�@U<�}����$�6�H�Z�
��^�^ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x�������������� ,>Pbt� ��#�����`(:L�2��P+�imih��0�A�B Ѓ�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?OO*O<ONOYG�w'cYO�O�O�O�O �O�O__&_8_J_\_@n_�_�_�_�_�Z�B��_�V�_i���A��_/m	12�345678�r�`!B  �
/h�@��jo|o�o �o�o�o�o�o�o q�O #5GYk}�� �������1� C�T�w��������� я�����+�=�O��a�s�����V�BH ��П�����*�<� N�`�r���������̯xޯ�[�;�j�� &�8�J�\�n������� ��ȿڿ����"�4�F�]�D�_wωϛϭ� ����������+�=� O�a�s߅ߗ�Z����� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1C�gy�� �����	-�?Qcu���U g`���`�//�mI"C��A�_J �  �qH2uB�gb%)
�Pdq#�
?`��R2��/�/�/,�/�+pM$ZO���/0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O?�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_��_�_ ooG!�$S�CR_GRP 1����� �t �G!� R%	 _Ra�Zb kbdd�f%f!�ekwgp�o�o�o(-�a ~�bD�` D��.�qcw�k<R-�2000iB/2�10F 5678�90� @tX� �RB21 OpC#�
V06.10 �zp�hKa�br#�u�vZa�fIa�cIa3Df!�ahj�a�y	�r��
��.�@�P����H��r�r^g��vN��`�pT@�q(à����0WB����,�5va= ���-�V>�ź�C4aBdX��@�H�P�  <���� @|�à�wZ`�OG!�o��o1�.'"��{h�p�Y
%���w`B���B� % ~�ǐ�vaAL ��G  @G ��va@�`ʟ  ?���v�: �򟨛vaF@ F�`�%��I�4�m� X�}�����ǯ��믖i ��������%�7�B�E�گ��v����� ӿ��п	���-��Q� <�u��/���c�o����Bi
����C#�@㑇�� ߘgΟ@�B��P�1234@Ns`׀h���C$A�g�Ra��㏛cd!2�rG! ���������2�>�P�� P�v�(|���� Ibp`�tZ`�}�{ yi��gϩo�i7��P�����7uIn�depe��nt _Axes Qs	�� ��n�f�w��s�w 3i��r���j|� ���c��	�vaC�s3/A�� Z��~iϢ�S�� /������/���F/ 藦�t/��/��/�/ �/�/?�/?=?(?a? P�:�p?�?�?Z��?R? O�?'OOKO6OoOZO lO�O�O�O�O�O���� #_f�����k_}_�_.�Rٺ_\�n�~�o�� L$o7o��boto�oUo �o�o�o�o�o��S�����_�� :��._��������� ������p�$6H Zߏ���'��� �o�~������Hoh ퟀ��#��G��h� 
/��./P/R/d/�� �0�1��U�@�e��� v�����ӿ�?�?��� ��?Q�Ŀu�`ϙτ� �Ϩ���������;� &�_�
�_m��F_X_ �����_�_�_�_�V�_w�o������o �������+�=��a�s���$6xBT�� ��3��W� ��,�>�P�b���� ������ΏSew� �:�L�^����// +/��ܟa/��/�/6� �/Z��/~� ?��įƯ دZ?|/�?�/�?�?�? �?�?�?�?#OOGO6�  �VOhOzO@��O8O�O �O_�O1__A_g_R_ �_v_�_�_�_~���_ L����Qocouo�2�8�J�8ff��o��4/ Z�Wi8y���������$�SEL_DEFA�ULT  ��_��P��MIPOWERFOL  6e.�7�oWFDO#� .���RVENT 1O����,��`�L!DUM_E�IP����j!?AF_INE"�Ə��T!FT����伏�!�>� ���e�!RPC_OMAINf�H��T����x�VIS��G�������!TP�P�U����d�I�!
�PMON_PROXYJ���e8�����c���f���!R?DM_SRV⯯�9gЯ-�!RZ�I����h�y�!
z�M䬯��ih�ſ!R�LSYNCƿ��8���!ROS̛�8��4 �]�!
�CE�MTCOMd^ϲ�kLϩ�!	r�OCONS�ϱ�l�� ��,�������B�g� .ߋ�R߯�v��ߚ��߀������?����R�VICE_KL �?%�� (%SVCPRG1r�D���2����3��D���4
����52�D7���6Z�_���7��D����8������9������D������' ����O����w��$� ���L����t���� ������?����g �����=���e ���/��//�� �W/��/��-�/ ��U�/��}�/�� w������B?�?�� �?�?�?�?�?�?�?O O?OQO<OuO`O�O�O �O�O�O�O�O__;_ &___J_�_n_�_�_�_ �_�_o�_%ooIo4o [oojo�o�o�o�o�o �o!E0iT �x�������M:_DEV ~���MC:�����%�~�L S  ���i��!��OUT�`�:�!�R�EC 1�d5L���   �j 	�  �݁ ���"���������􍶃 �� ���� ��4�C�
 �W
O6 ���� �U� �� �s�t_d5T������.�b �  �瑁�7�U� �7��M�x ��$M�p��	h�����UM�����<��љXQ� ]�x�����B����XD�џ�\M�?���)���o7�� ��M�) �e �U� U"i�� ���L7���}�RW9�]��* �v �� � �{�U}� ����� �iJ �m!���� �U27��M�� �g ��Hٯ	� ��7������M�Đ �.��kw]��M��q�f=� �� ��)� *t�t �zI��Q����a��7��M��7���7�孿�a����q���7�*����#�����r�@�]�P�!j �Ȱ ��q��� E!n �u�6�������Ϳ߶)��p���7�.��1\f�����]�� �)P �ȑ �͡1ϫ * ���+ �cB �^���!��� ���7�3���D� ��-�Sy@�(Ѽȁ���!\-�K�ݚ�dͣ������b��yɟۖ����Y�M�<�u7���ٯU�I0]��Ť��ѕ��� ���Ť= ����)ߪߒGM������Z� �]���V7�_�6�)�p�U���� �
T��C��  �� V�Y �� ��]�+��7��7��M����M�d	���7�/�E�7���D�v��WB��]�� �l ���B �'Ł�|�!���K��1�o��ߒE� ��7���������7�6���V�R'-7i]�ȑ� �쐔�|ѵ�� �ȡ}BI��UϷ���pɹ}�f����������_�������A	/Q'�]��M�`�e] �� �$� �A �w������gyd����������� ������) Q-]�\m�X �� ��� ��� F��iB6��#5���Y��� ������
�(^��СPѣj �� �ə I}��u��������*鰀������ ��^cQ(r�a���p �<!��D/  > � �������l/~/�/�U鰤���7�� Z���+;�]��M�U
 �[ �� ��ɡ �/��["���?'?�9?�`����|����� � ��9P�+��]�� �� ���� wy�����k��Ń� �1����ß՜ ���~�C�z�J7��J�Kd�]�~
� ��q��B�O ��|�H����?��?�?�D����#�� � �����IM!C\�������� �U��O C� �{6� �rE_k�A_��鰜������� ���ឡYNoE]� ��J �A �| � ���_ C�@A�AL�,��_._@_hⳠ\ � �� V���+��D� ���o���1/S�F��O�f�6r[",��Mi���T����ak����/P)�}{�JA���e����O�����K�]� ����ý��������"j`��	�g����i�0G�Y�ß���ş˟ ����ϋ��m�ז�ڕ�[���sT[�����o�J񯫯���R��#��k�NVN��+S�Z��W������+!ɿϿ���N�N���.����	��s�1���]ϻ�5�OJ��T6 �Iw(���ϣϵ�����`!�'��o���@q�O�a�����$*�߷�����W�E� {�i�����ɯۯ�� ������S��w�Y� ������������� +O=_as�x��wCL�Lm�+Ajg�)Ӛ�1x7!Jׅ#���&�ϫe��� ���+/�;/=/O/ �/s/�/�/�/#�5�? /??G�9?#?�?� ���?q?�?ٿ�?�?O 5O�/YOGO}OkO�O�O �O�O�dL_H)__ M_8_q_�_6��O�_�_ �_�_�_�_"o4ooXo Fodojo|o�o�o�o�o �o�o0TB` �l������ �,�>� �b�P���t� ����������� :�(�^�L�����v��� ��ܟʟ�� �6�� F�H�Z���~�����د �̯���2� �B�D� V���n���¿���Կ 
���.��O�_,�v�d� �ψϾϬ�������� �$�*�<�r�`ߖ�x� ���ߺ������� � J�,�n�\�~����� ��������"��F�4� j�X�z����������� ����BT6x f������� P>tb� ������// /L/./@/�/p/�/�/ �/�/�/D�n_'??K? 6?o?Z?�?�_X��/ ? �?�?�? OODOVO8O zOhO�O�O�O�O�O�O �O�O.__R_@_v_d_ �_�_�_�_�_�_�_�_ *ooNo0oBo�oro�o �o�o�o�o�o& 68J�n��� ����"��2�X� :�d�j�|�����֏ď ����0��T�B�`� f�x���������ҟ� ��,��P�Fϸ?^�`� �������ί���� :�(�^�L�n�p����� �����ܿ� �6�$� Z�l�Nϐ�~ϜϢϴ� ��������D�2�h� Vߌ�zߘ��ߤ����� ����
�@�.�d�v�X� ������������ ��$�*�<�r�`����� ����������  &8nP~������f��$S�ERV_RV 1-�	8��0(	\ �n���!3�TOP10 1��=
 6 ��02 2�0 r�0 s�06���0 �0�6 &2" ���06r _"$�E�YPE  �1�H�01�HELL_CFG� �t&�0�?�X"�/�/ %RSR�/�/�/??:?%? ^?I?�?m??�?�?�? �? O�?$O5MDD<I�; �E%5OvO�OCE?M� �O�B�@K�D\D!d�O�"�)]!�#HK 1�+ �O<_7_ I_[_�__�_�_�_�_ �_�_oo!o3o\oWo�io{oC}&OMM ��/�o|"FTOV_ENBi$Et*�OW_REG_U�I�o{"IMWAI�T�b�I{OUTrvDyTIMuw��WVAL,>s_UNIT�c�v�t%]!LCpTRY�wt%1MB_HDDN 2�k )P��� ��>�5�G�t�k�}�𪏡�̌�qON_ALIAS ?e�iLhep���(� :�L�D��w������� X�џ�����ğ=� O�a�s���0�����ͯ ߯񯜯�'�9�K��� \���������b�ۿ� ���#�οG�Y�k�}� ��:ϳ��������Ϧ� �1�C�U� �yߋߝ� ����l�����	��-� ��Q�c�u���D�� ��������)�;�M� _�
�����������v� ��%7��[m ��N���� �!3EWi� ������// //A/�e/w/�/�/F/ �/�/�/�/?�/+?=? O?a?s??�?�?�?�? �?�?OO'O9OKO�? oO�O�O�OPO�O�O�O �O_�O5_G_Y_k_}_ (_�_�_�_�_�_�_o o1oCo�_Toyo�o�o �oZo�o�o�o	�o ?Qcu�2�� �����)�;�M� �q���������d�ݏ����%�Ѓ�$S�MON_DEFP�RO ����N� �*SYSTEM�*Ё�>�REC�ALL ?}N� ( �}׏����ԟ��� ���/� A�S�e�w�
������� ѯ������+�=�O� a�s��������Ϳ߿ 񿄿�'�9�K�]�o� ϓϥϷ������π� �#�5�G�Y�k��Ϗ� �߳�������|���� 1�C�U�g�y���� ����������-�?� Q�c�u���������� ������);M_ q������ �%7I[m  ������~/ !/3/E/W/i/�z/�/ �/�/�/�/�/�/?/? A?S?e?w?
?�?�?�? �?�?�?�?O+O=OOO aOsOO�O�O�O�O�O �O�O_'_9_K_]_o_ _�_�_�_�_�_�_�_ o#o5oGoYoko�_�o �o�o�o�o�o|o�o 1CUgy�� ������-�?� Q�c�u��������Ϗ �󏆏�)�;�M�_� q��������˟ݟ� ���%�7�I�[�m� � ������ǯٯ�~�� !�3�E�W�i���z��� ��ÿտ������/� A�S�e�w�
ϛϭϿ� �����ψ��+�=�O��a�s���$SNP�X_ASG 1��������� P 0 �'%R[1]�@1.1z� �?�r�%����<�Q����_*_�G��Ƕo�6�w� �.�f��֦����� �ǯ�#����� q���7��$�E&�g���KV����ǟ8����֡0q������!�0��'� t�W���� �� �8v��/�����v��
�12G
̈́6w����� ׆1��� �lG�/�����6/ �Qq�&/g/�Q<V/��/�����/h	��/�/ ��/&? ׄ#��?W?I�F?�?��&�v?�?�2�Y�?�?��ϴ�?O�׋OGO����6OwO��?�OY�|x�O�O��	�O_�n�qM�O7_��	�&_�g_��߅/�_ �Jc�\�_�_��5O��_ ��u?&o��51OoWo�O�Eo�o� �]o�vo�o��1��o�o�zb��� �ޒ%/F יC�Ov����f�:#� ��7�/�� �����7��'A1J&�g�ֵ���� ע�%��Ǐւ�A/������4�8�'��~j�W���@��� ��I1�v�����>w����ZwN�֟��R�8u�F� ����6�w�ƪ'�f���֑�1���ׯ��6�O�F א��6��I|&�g� �'���ߋ�̿�Ѹ����� ���'Ϫ��]���#1tFχ�և��R���PARAM ������ �	B�P<�P!�I�D����OFT_KB_CFG  ]��ԉ��OPIN_SIM  ����=�O��a�Q ��RVQST_P_DSB&�������h��SR ��)� � & �FOLGE125� .����0021�A��Ī�THI_C�HANGE  �E��GRP�NUM� �O�P_ON_ERR���I�PTN �)��C��RING_PRt1�U���VDT+�' 1�ɑ@�@�� �F��������� �1� C�U�g�y��������� ������	-?Q cu������ �);M_r �������/ /%/8/I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_P_a_ s_�_�_�_�_�_�_�_ oo'o9oKo]ooo�o �o�o�o�o�o�o�o #5GYk}�� �������1� C�U�h�y��������� ӏ���	��.�?�Q��c�u�����e�VPRG_COUNT���|��ƒENBđ���M�4���UP�D 1���T  
����B�T�f��� ������ׯү���� �,�>�g�b�t����� ����ο�����?� :�L�^χςϔϦ��� ��������$�6�_� Z�l�~ߧߢߴ����� �����7�2�D�V�� z������������ 
��.�W�R�d�v��� ������������/ *<Nwr��� ���&O J\n����������_CTRL/_NUMГ!��!"GUN%" 2}�0��  1$(4!!4!/s$
1$Ւ(#�'�/�/�/�/�ÐYSDEBUG�А1�� d�� S�P_PASSЕ�B?;LOG ��0�� �J1�^��k$[=��%UD1:\x04.12_MPC6?� c(�?g=x82��?�2SAV �9=�!n%&x8S�V�;TEM_TI�ME 1�R+ �( A4"0靟&~I��! gG��sHEO�O{@�:�O�O�O �T1SeVG S+�ѕ'���PASK_OPTIONА0��ߑ'Q_DI0�ߔ�TBCCFG ��R+�=�.�_`�_���!�_�_�_o �_5o oYoDo}oho�o �o�o�o�o�o�o
 C.@yd��� ���	���G�6� �i�{��X�����Տ �����0��=P�!� G�5�k�Y���}����� ßşן���1��U� C�y�g�������ӯ�� ����	�+�-�?�u� [�F�������˿ݿ[� ���7�%�[�m�� Mϣϑ��ϵ������� ���E�3�i�Wߍ�{� �ߟ����������/� �S�A�c�e�w��� ������+�=��� a�O�q����������� ����'K9[ ]o������ �!G5kY� }�����/� 1/��I/[/y/�/�// �/�/�/�/�/?-??? ?c?Q?�?u?�?�?�? �?�?O�?)OOMO;O qO_O�O�O�O�O�O�O �O__#_%_7_m_[_ �_G/�_�_�_�_�_{_ !oo1oWoEo{o�o�o mo�o�o�o�o�o /eS�w�� �����+��O� =�s�a�������͏�� �_	��9�K�]�ۏ ��o�������۟��� ͟#��G�5�k�Y�{� }���ů���ׯ��� 1��A�g�U���y��� ��ӿ������-�� Q��i�{ϙϫϽ�;� ��������;�M�_� -߃�qߧߕ��߹��� ����%��I�7�m�[� ������������ ��3�!�C�E�W���{� ��g��������� A/Qwe��� ��$TBCSG_�GRP 2����  ���  
 ?˃�@����  <N8r\� ������� /,//P/:/t/�/l/ �/�/�/�/�/?�/(? :?$?^?D?n?�?~?�? �?�?�?�?O�?6OHM�A��*SYST�EM*� V8.2�306 qC4/2�x@014 A �t  _F_GF��� PARAM_T�   �$�MC_MAX_T�RQ��$�D_MkGN�CC� AV�I�STAL�IBRK��INOLD�FSH�ORTMO_LI�M	Z�M�EJPTP�L1CU2CU3CU4�CU5CU6CU7CU8��A `�A��A�� �_AC�CEJR�WTQ�SP�ATH�W�Q�S�Q_RATIO�B�S�@� 2  	$C�NT_SCALEn	ZSCL�CIN�Q�_UCA��bC�AT_UM%hYC_ID 	*cB`_EKPGjTPGj]P~G`PAYLOAW�J2L_UPR_7ANG�fLW�k�a��i�a�ER_F2LoSHRT�gLO�d�a�g)c�g)cACRL_Shpgzd�B�HVA`  �$H�B:rFLEX�7s�@Jb�@� :$aLE�NKQguTQ$DEjx�t|s�R�X�p�z�SLOW_AXI^q$F1aI�s�2�x1�q�u�wMO�VE_TIMd_?INERTI%`:p�	$D	�TORQCUE�Q!��p�IHPACEMN�`��P�s�E^�V�p�A/�8x�@�x�TCV���@@��A�������@T.��@��J�A�����M	�(a�(`J_�MODa�p� �R�@�gq2�@P��^�Eo�0`J��X�p�A�RU�?�JKh.�����KKSVKTS;VK]SJJ0�KS�JJTSJJ]SAA6KSAATSAA
�fS3AAoS�AN1ǌ<�𒋳@�@PE_NU�QΈVqCFG��A � $GoROUP�@SK&c�B_CONFLI�C�dB_REQUgIRE.q�qBU s_UPDAT�v� �ELk�� Τ�$TJ�P�J�E�@CTRa�qT�N	�F˦��HAN�D_VB8rVqO�P�U $]�F2��F
�TSCOMP_;SW&a  $�@�F� $$M�`�IR�C|��A��x��LR��A_}b�FDļ��MA�LA�LA�KA� [Ұ�KD�LD�KD� [P�PGR�Gp�S�T�Gp��Ip�NXDY�`R�@�E��ڵ�`  `�g�q�g�a�g0�<Q@��p��UPKUTU]U`fUoUxU�U�R$�Vr��T r�Wt�R �%�n�TPy�ASYIM�U:p� �V�P8m�ao_SHo�g 4d]��C�>oPoboto�cJ�l>P�j^�T�i.
�_VI&����>��V_UNI�c��TS�aJ��������l ���e����m�y>P�1a���GtOs���|�TCPPI�R�A  ��EN�ABL�p����$TCDELAYݱ�g�t��SPEE�4P  X ���I�N� ސ��� �GP����Q���q�@M}PڢPROG_��N�YPEڡ��_z��	 |�m���SE� s��m���' ǦWA7RNI��EN&����OTF�qj��_TL���MAARSCW���SPDz�
 �������EARTBE���ET��z��ӝPPARGAT��F�LG�u�|sS�@E
�@R&�6�%�a8os6REAJVX�TR�� OUT�AC p렜��� E�̢�ID`�(d^�Uc�A�`��޵��G�Q# �PH����<��{I�$D=O� ���z�� ��I��A ��J �p��W#�۠�L��q�� �[ T�MES���R���T P��"@Pl���#��(�!�)T"�m� $�DUMMY1]Qo$PS_�pRF�p�g@$�&��FL�A|��2�GLB_Tu�k*5���()���8!�����Q�STT��SBR��PM21_V�T�$SV_ER�`O��p3�3CLD0p2A�^����GL��EWΦA 4��$��$ZݲW�3���`rP�As %b  ̳3]U�5 ]�N�0��$GI�}=$�1 / �1�0�A L��F�W}$F�EFN� �M�NcF]IJ�TA�NCb L�J� RǱ +!$JOINT�����1M� �Q��FECE�q��S�b��*B����Q� �pU�S�?��LOCK�_FO�`[�� BG[LV��GLXT  �_XM`�AEMP��@�� -PB2�@$#US�!�0p2*��4�QQRW��@QQ�S�CEj�CrP $K���M#TPDRqA�0�T�AVEClp��V�@IUQQVQH=E�@TOOL�s�S�V�tRE�PIS3�|s�T64�)`ACH4� ���QON��$�29�"�PI� � @$RAIL_�BOXE���R�OBO"T?�r1H�OWc>d� aROLM�"ge_�
dxb���/`�p6�O_F��!   �2�Q^q]�Ot�R�PO]r!�b�p�A�`��1~X2MU�֡��,�@	 IP#VNK��R�/b�Q
�QQ�`�PCORDED�@���`�1���OY   D )0OB�٣�@�dwSq�#E Sr�ۡS;YSSqADR =Q�TCH��  �, �A�A_D��th�*�@TPVW�VA�� � ��P�2kPREV_�RT��$EDI}T�VSHWR�����$�K��IND�� `;�$��D�&�[�U�6��KEp��� �l�JMPpp�Lj@�TRACUE)[p�I,P5SڢC �NE�Pۡ���TICK�S��M�o���HNR1� @]p��L	_G8K&f��STY�aLOD1����~�_ t 

 G�uS%$�qD=� SFp!$��8��!�F r�P��LSQU�aLO���TER�C� ��TSz� @h0�� p���㡼Q,�O� �#dI�Z4A��! Cx�"!�oUTPU���1�_DObB�pXS:�@KjAXIP��c�VQUR���0i#$ATH`�~vK���_�P�rET��P Rlp��%O�F��P�A������$ cc>  �-"SR3� l ѐu��A�������� ����ù�ӹR��� R��R��d�~�B�d�H���҂�C翐�C���� �2�D��SSC�,0 ! h�0D�S�� X}�AT���<�� ~���"AD�DRES�SB�S�HIF�HP_2C�H� zqIK0���TXSCREEUr�"	 k�TINA�3@��D-!����T0# T���0'Ҁg00�^��r^��RROR_vA��(�h$v�AUE5$$ ����q0S�1�qRSM<��T�UNEX��j���S_�3��G������G�C�B���? 1# 
z���%="�2��MTJ!�Lv�m�w0O�D���UI_� H>P� & 8e�w@!_T���f� R���BXcg�"@R�O���T0'���7$B�UTT��R RraL�UM��u���ERV��R�Pa@��S1(z{ ƠGEUR&SiF���A)� LP���E��C�)#�S�1�Pc�1��P0�5.�6.�7.�8����a@P���%�Q�AS��'R�USR�4') <Z0� UB�A9I΀@FOC�Q@PRIΡm`�� �TRIP�m�SUN$ 5$*	@t�0$ kcj��HR����� +a��� �G� \��1���\O	S�qR��V�H�QS1,�?�3�>���`HRU�S1-����8��HOFF!PT0�.[p�O' �1,�09-�0G�UN_WIDTH|�B�B_SUB�"�p0�SRT� �/0��vA�` �OR`�'RAU��T�����VCC�М�0 ��aC36MFB�124�AVC/0.D1�h %bTq�� �4.��c)�C�`	%�DRIV���_�Vu�,$(��@D��MY_UBY��$V� vA�� B�tC�#�QtB�i0pp+��"L7�BMv�1$��DEY!��EXG�n��Q_MU��X�10orbҲ�}GðPACIN΁}�RGC�52�20�32���!RE{�����Q�B��2�02^�TARG�@P1R�c0�`�R� �03 9d��_�FLA΀r�	�"N�RE�#SW0_A1�@�@�!��O���A���3�E���UB�a�@�hV�HKG�4���:`����05�!CEA���+GWOR!P�5 ���MRCV�5 U���OS�M!PC2S�	hB`3hBREF F�FqF\A�0�࿣�0 ��mJ�A~J�A�K�EqFO_RC,KXEKV�S���']#�OB���6 �$���1؄8��b%�pROU�[2<�# 1z52��2�P$���� �΀�3��2���Kq�SU�L��4;r��� 5� �P@�3�cN�f ��f��c�PL�#5e`�#5e��Ag���$>��70 &��ǡ�4� ��C�`+�LO �A�d�a� �iu��`ܓmC�pMI��FR�hqTj��fR[$HOh�z�r�`COMM'#��OB�v{X����؇VP]2�Hq_S�Z3cQu6/cQu1�2��Nx0Lx�`LxW�A�eMP�zFAIj�`GT�`AD�y��!IMRE~T�r_��GP��� ��&A�SYNBUF�&V�RTD���qσOML��D_�:�W��P�ETU�#�`Q��0�ECCUP8V�EM:0�e���gVI�RC�q2�le�8|u��0CKLAS^?	�VLEX��%9/�����	��LDLDE�FI@<� �r���S@��TpT�Q��:����T�1�'�����V�� ;`��L����{,�"UR�3�0_R �p󔟑�!���U3�/ �/�$�`7���0Ғ �sTI�Q��SCO�� �Cz�4;#6;� ;�;!�;/�//%*ᢕ���D�SЧ@� f0SM�<)���J*��%���q�=)G�eL�IN���W�@X9SGAq�>  ��N��BPK�cH��HOL��� S@ZABCB}?v2`�XS�@
�_ZMPCF}@<�d��2��l!LNI�Ƙ@
L��� ~A ����q+@��CMC�M0CKsCART�_ٱ�DP_�� $J����������S��S��BUX9W� ��UXE�!A�<��9��d�J�\ɴJ�l� ��ZPץBc ��b�`��uY!�D" Ca�:���IGH&3G��?(!�!��A�T|���D � T�,�A~�$B�PK�'3PcK_a�	c�RV�`qF��Ba�OVCYЀ���TU�O0��j�
�RI��1uD��TRACEx�V
1^�͐�PHER��E �,!������ɸ�$�Tb� 2������ d ���? �	 HD�)ˀ� (�CX��0�)�(�$�BE��O�Z�$�33]3x���<�|Z�8\�&�8��.�����C��� CA��C0�������tP�P��#�2�6���sz����K���@����� ������&C n��p��	�V3.00�	�rb21�	*�� ����
fffjtW�^p	 ��   ?���Cz�_f�x�� �� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?O��	 O2OO ^OlI0pO�ODlO�O �Kz�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>PbO>O �JO���O��O� (��O0�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯t� ��.��B��v�舿���J�� v��  f+���2f�G����	2 ?�*�c�Nχ�rϫϖ� ���������)��M� 8�q�\�nߧߒ��߶� �������#�I�4�m�@X��|�������� ������8�#�\�G� ��k������������� ��"XC|� ��I�s����� !E3UWi� �������/ A///e/S/�/w/�/�/ �/�/�/?�/+??O? a?k��p?�?�?>?�? �?�?�?�?OOBO0O fOxO�O�OZO�O�O�O �O�O_,_>_�O
_t_ b_�_�_�_�_�_�_�_ oo:o(o^oLo�opo �o�o�o�o�o �o$ H6X~l�� �����?�&��? �h�V���z������� �ԏ
��.����d� R���v�����П⟜� �����*�`�N��� r�����̯��ܯ�� &��J�8�n�\�~��� ��ȿ���ڿ���4� "�D�j�Xώ��:��� ��tϢ�����0��T� B�x�fߜ߮����ߐ� �������P�b�t� ��@���������� ���L�:�p�^��� ������������  6$ZHjl~� ����� 2�� J\n���� ���/
/@/R/d/ v/4/�/�/�/�/�/�/ ??�/<?*?L?r?`? �?�?�?�?�?�?�?�? O8O&O\OJO�OnO�O �O�O�O�O�O�O"__ F_4_V_X_j_�_�_�_ �_p�_ o�_�_Bo0o foTo�oxo�o�o�o�o �o�o,<bP ����v��� �(��8�^�L���p� ����ʏ��ڏ܏�$� �H�6�l�Z���~��� Ɵ���؟���2� � B�h�o������N�ԯ ¯����.��R�@� v�������j�п���� ��*�<�N��^�`� rϨϖ��Ϻ������ �$�J�8�n�\ߒ߀� �ߤ����������4� "�X�F�|�j���� ���������$�6��� V�x�f����������� ����,>��NP�b����  � � �����$TBJOP_�GRP 2W���� ?���C�	�E�� ������X��y�^� �,X�� @� ?����D)̴C2
C랔���wB;�(����;S��!���<p�S�>�+�L?%H�?$+�LB�g"B:��'/2'���j/�|%<?D!?���?L�#C  B�Z'�/:/L/^/܀/4CX�2)��;�ŗ-C?�~B��~�/Q?�Cd6����C�p"�*tP���6�?�'�;����CA�?=���?p��1Cu�CP�R?�?d?�v?�6h4O�6;��?)�2 ?W^��PAC;֭C���?qO�?O B�E�O�7Kl��2333�?fff?Y-Z�@rO�O�;�%_�' 4__,_Z_�_f_ _�_ �_�_�_�_o�_�_:o@To>oLozo�o~D����� ��%	V3�.001rb21�*�`���w F�� �F�. G
� �G(� GG� �Ggs G�� �G�v G�^ �G���G�@��G�; G쑀�G�C�H	(��H� H���H&��H1��H;y� r?� �FM4 Fj0 �F�` F�v �F�V F� �G> G7� �GZj G�l �G���G����G�� G�� �G���HS@�H��H0) �HB�@=� <���l?� W� _�@j����
�?�  ��oK�y� `�\�n����G����ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤߪ y���߬߮  !p���(�:���^�p� �����	����� �j�)�����u�?� ���������������� ��);M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?OO+O=OOOaO sO�O���߳O��S��O __�O�OK_]_o_�_ �_�_��_����_1� Y�#og�y�ko}o�o�o �o�o�o�o�o1 CUgy���� ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W�i��O�O���O 7_տ�����Ϳ/�A� S�e�wω��_���_�_������$TCPP�ACTSW  �e���I�R e����CH%�SPEED 2�� C�e�  ��ͮ��_CFG K	2�?Ѵ����!Ӯ��_SPD��
�>�  ֽQ?�:�o��p�������NUM������
��OUT ;2��
  ���� t��n������� ������/�"�S�F�X�xj�|��ZERO���  ���ESTPARS�?�����HR��ABLE K1���Ҋ���*���������Ѫ����	��
��P���������4���RDI��<��&8J\�O ����0��	S��� �
�// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?�����z�w� ��Yk}���X��n2/� 2�P`��0 3�4�����2�A@��`�IMEBF_TT��p�5�զ�CVER2��!ѯF�ќ@R 1��8ﴰ֌	] 	a��7a�6�����OR�P�P\�$_hY��KuPU�0[�\_�[QR[Ĕ_�_�_c��_�_�_�o�Gh�S�
��H[Ǭ�DooXY�<oNi��\`�`o��to�h�ި7) �o��oEB�oVˬo�
;S�T��inX}�H�i�]��~�n�rV����S_E�bV�4��oX��l��~���Ҥ���d��V�܏F�T_�������93�3�E���c�h�z���� }��������������u?��"���_[8/�Y�k�'���������*B��ί���#������g�9��K���`�r�L��w������D.�!�@��� �MI_CH�AN�G 
�DBG�LVL�G���E�THERAD ?���i����0�r�:eu�4:37:14:f0 r�Q1��5���3P�RP�6�@!��!�������SNMASK�^���o�255.$�0��#�5�G߁��OOLOFS_D�I���L�ORQC?TRL �ɦ3�:��5�T������ ��0�B�T�f�x�� ���������������;�*�_���PE_DETAI<ȉָA�PGL_CONF�IG WIgA��?/cell/�$CID$/grp1c�?�c�����(�����2(]@o���4��3����)���4 0ew���<�� ���/ /2/�V/ h/z/�/�/�/?/�/�/ �/
??.?�/�/d?v?@�?�?�?�?���}S?��?OO*O<ONO  O�uOTN�R?�O�O �O�O�O_L?)_;_M_ __q_�__�_�_�_�_ �_oo�_7oIo[omo o�o o�o�o�o�o�o �o3EWi{� �.������ �A�S�e�w�����*� ��я�����+��� O�a�s�������8�͟ ߟ���'���K�]��o������������User Vi�ew ��}}12�34567890 �����0�B�J�Ӱ��j���ΩK	�?�� ��Ͽ��� e�w� բ�	��_�qσϕϧ� ���*ψ�SN��%߀7�I�[�m����ψ�5 �ϼ���������u�7�}�6��p���� ����)���}�7_�$� 6�H�Z�l�~����}�8������� 2���SY lCamera٪ ���������BE�.@�Zl`~�����  r ���//(/:/L/^/ �/�/�/��/�/�/ ??$?K�rBɻ/ p?�?�?�?�?�?q/�?  OO]?6OHOZOlO~O �O7?I7��'O�O�O _ _$_6_�?Z_l_~_�O �_�_�_�_�_�_�OI7 ��_Jo\ono�o�o�o K_�o�o�o7o"4 FXjos^��o� ������o2�D� V��z�������ԏ {I7�k� �2�D�V� h�z�!������� ��
��.�@��I7�� ן������¯ԯ母� 
��.�y�R�d�v�������S�e�98���� �#�5�G��X�}Ϗ� 6�������������
��	t0��Z�l�~� �ߢߴ�[������ߣ�  �2�D�V�h�z�!�3� y {�������	�� -���Q�c�u������ ����������t��� ?Qcu��@�� ��,);M _@�S;���� ��/�)/;/M/� q/�/�/�/�/�/r� �Kb/?)?;?M?_?q? /�?�?�??�?�?O O%O7O�/�+k�?�O �O�O�O�O�O�?__ %_pOI_[_m__�_�_ JO��{:_�_oo%o 7oIo�Omoo�o�_�o��o�o�o�o�]  �Y>Pbt��������� �  y?���B� *��]>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D�pV�h�z�(x  
�`�(  �2p( 	 �������ο ��(��8�:�LςϠpϦϔ��ϐ�z �^o�!�3ߦoW� i�{ߍߟ߱߸S���� ����F�#�5�G�Y�k� }��ߡ��������� ��1�C���g�y��� �����������	P� b�?Qc����� ���()p M_q����� ��6/%/7/I/[/ m/���/�/�//�/ �/?!?3?E?�/i?{? �?�/�?�?�?�?�?O R?/OAOSO�?wO�O�O �O�O�OO*O__+_ rOO_a_s_�_�_�_�O �_�_�_8_o'o9oKo ]ooo�_�o�o�o�_�o �o�o#5|o�ok }��o����� �T1�C�U��y��� ������ӏ���	�� b�?�Q�c�u���������@ ��ȟڟ������)f�rh:\tpgl�\robots\r2000ix&��b_210f.xml��P�b�t����������ί���� >�dummy"�;� ?�Q�c�u��������� Ͽ��
��.�;�M� _�qσϕϧϹ����� ����*�7�I�[�m� ߑߣߵ������������)�;�M�_�q� ������������� �%�7�I�[�m���� ������������! 3EWi{��� �����/A Sew�����t��;� ��88�?� �"/�/@/B/T/v/ �/�/�/�/�/�/?�/ ?B?,?N?x?b?�?�?��;�$TPGL_�OUTPUT ���  ?O���3;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_@m__�_�_�3 �@�2345678901�_�_�_�_o o (c��_Ooaoso�o�o �oAo�o�o�o'�j}1Yk}�� 9K�����1� �?�g�y�������G� �����	��-�ŏ׏ c�u���������U�˟ ���)�;�ӟI�q� ��������Q�c��� �%�7�I��W���� ����ǿ_�տ���!� 3�E�ݿ�{ύϟϱ� ����m�����/�A� S���a߉ߛ߭߿���i�A}!��+�=�O�a�r�@/���* ( 	 �_ �������%��I�7� Y�[�m����������� ����E3iW �{������/�V� "7e wS������R P
//�@/R/0/v/ �/��/�/`/�/�/�/ �/*?<?�/`?r??�? �?�?�?�?H?�?O�? OJO\O:O�O�O�?�O �OjO�O�O�O"_4_�O  _j_|__�_�_�_�_ �_R_oo�_BoTo2o do�o�_o�o�oto�o �o,>�obt �����J\� (��L�^�<������ ��ʏl�ڏ �ޏ��6� H���l�~� ������� ؟�T��� ��V� h�F������¯ԯv� ��
��.�@���,�v� ��*��������������$TPOFF_�LIM K|�ӱ��|��Nw_SV�  x��%� �P_MOoN CG��*�|�2x��STRTCHK C�E��M�VTCO�MPAT:���I�VWVAR Z�Y��h��� ���|�m��_DE�FPROG %���%FOLGE�12��Y�t�_DISPLAY���/��INST_MSK�  �� k�I�NUSER��q�L�CK�܊�QUIC�KMEN��q�SC�RE�C��tpscq���!�h&�%�7�_;�ST���E�RACE_CF�G Z�����	�
?���H_NL 2��#���� ���������"�4�F�X�j���IT�EM 2�� ��%$12345�67890���� � =<�������� G !����� Jӫ�k���� �);_�/ U����	� 7�	//?/�� �A/��/�/�/3/�/ W/i/{/�/M?�/q?�? �/�???�?A?Oe? %O7O�?MO�?O�O�? �OO�O�O�OaO	_�O �O�O#_�Oy_�_�__ �_9_K_]_�_�_�_So eo�_qo�_�_�o#o�o Go}o/�o�o| �o��o��SCU g����[����� ����-�?���c�� 5�G���S�Ϗ��w� ş)����_������ ^���y�ݟ�����ů 7����m�-���=�c� u�ٯ�����!���E� ��)ύ�Mϱ�ÿտ Y�q������A���e� w�@ߛ�[߿�ߑ��Ϡ���+��߀�S��|��F��  u��F� ��P�F�
 �]��j��(�UoD1:\������R_GRP 1 ���� 	 @P������1��U�C�y�g�������s�����������?�  )I7m[ ��������3!WEg�	�ա�q��m�/ �'//7/]/���/�� �/���/�k�/#? ?G?5?k?Y?�?}?�? �?�?�?�?O�?1OO AO���O��Oe/�O �O�O	_�O-_k/Q_�/ x_�/u_�_QO�_MO�_ �_oo'oMo;oqo_o �o�o�o�o�o�o�o 7uOSe#_�_ ������M_3� �_Z��_~��_���� ՏÏ�����A�/� Q�S�e���������㟀џ�Eo5�G��S�CB 2!� ����������ϯ�������X_SCREEN 1"���
 �}ipn�l/X�gen.htm$�w����������P�Panel� setupü}�	index.STMÿ��1�C�U��̷
Robot ?Info e�9���ϱ���������  �τ�1�C�U�g�yߋ� ߯�&�������	�� -�߶�c�u���� ��4�b�X���)�;� M�_����������� ����x���7I[ m�6,����!3�W3�U�ALRM_MSG� ?D��Q�  RD������ /
//:/@/q/d/�/��/�/mSEV  �{�&kEC�FG $e�  �D7�A1   �Bȗ� Q�0��42B-��W;�$N246A�ڐ�WqK�28i2@�?��O��b?t2��z?t0 �=B�A<O_	2>.@O}z�J=�B2fpP=<��J>���T�f��>)��U:��~�!GRP 2%e�� 0N��:?��!�BPR;����@I>??G=ԎQ�,�0!�C��/�Om��O�O��O�OiI_DEF�PROw+F� �(%UP031� .%_-T0071�  %MAKRGO05<AQ_D%�/ _j_�_�_�_�_�_�_�o!ooEo�GINU?SER  ]�O�NoI_MENHI�ST 1&e�  �( P���./SOFTPA�RT/GENLI�NK?curre�nt=editp�age,FOLG?E020,1�q�o0*D�(�o�e�menu�b935,BPq���6HZ~153n��'�d9��p'�Z~74����������K�]��a37u�
��.�@����81��2m����D��F�-X��o�a1��5ȟ�,�>�I��o���4,8�����¯D�6a�a6o��� � 2�D�V�Y�므����� ��ȿڿi����"�4� F�X��|ώϠϲ��� ��e�w���0�B�T� f��ϊߜ߮������� s���,�>�P�b��� ����������ݯ �(�:�L�^�p����� ���������� ��$ 6HZl~�� �����2D Vhz���� ��
/�./@/R/d/ v/�/�/)/�/�/�/�/ ??�<?N?`?r?�? �?�?�/�?�?�?OO &O�?JO\OnO�O�O�O 3O�O�O�O�O_"_4_ �OX_j_|_�_�_�_A_ �_�_�_oo0o�_To foxo�o�o�o�oOo�o �o,>)?�ot ������o�� �(�:�L��p����� ����ʏY�k� ��$� 6�H�Z��~������� Ɵ؟g���� �2�D� V����������¯ԯ �u�
��.�@�R�d��Oz�$UI_PA�NEDATA 1�(������  	�}�/frh/cg�tp/respo�1.stm?_B�USY=TRUE� Save&AC�TION=101&C2=3p������  )pri9m�<�  }?�c�`uχϙϫϽ� )�� �������+�=�$�a� H߅ߗ�~߻ߢ���������Lv�� �    ��MĨ�vagmn�� *�m�������ual����O�  ��$�6�H�Z��~� e������������� ��2V=z�s�#� �������� ,>P�t�� ������Y/ (//L/3/p/�/i/�/ �/�/�/�/ ?�/$?? H?Z?���?�?�?�? �?�?=?O�2ODOVO hOzO�O�OO�O�O�O �O
___@_'_d_v_ ]_�_�_�_�_�_�_g? y?*o<oNo`oro�o�_ �o�o-O�o�o& 8�o\C��y� ������4�F� -�j�Q���oo�o֏ �����0���T��o x���������ҟ9��� ��,��P�b�I��� m�����ί�ǯ�� (�:�����p������� ��ʿ��a��$�6� H�Z�l�~�忢ω��� �������� ��D�V� =�z�aߞ߰ߗ���G� Y�
��.�@�R�d�� ���Ͼ�������� ��<�#�`�r�Y��� }�����������&�J1n����}������ ) �7��&cu�� ��$��/�� ;/"/_/F/�/�/|/�/ �/�/�/�/?��������$UI_POSTYPE  ���� 	 ��?��E2QUI�CKMEN  �T;c7�?�8RESTORE 1)���m0��?���?�3�?��m ODOVOhOzO�O/O�O �O�O�O�O�O_._@_ R_d_Oq_�_�__�_ �_�_oo�_<oNo`o ro�o�o9o�o�o�o�o �_!3�on� ���Y���� "��F�X�j�|���9 C�����1����0� B�T���x��������� c������,�׏9� K�]�ϟ������ί� ����(�:�L�^�����������ʿ�7SC�RE�0?�=�u1sc�0uU2�3�4�5ĕ6�7�8�E2U�SER����ksT�f�3f�4f�5fĕ6f�7f�8f�E0N�DO_CFG �*T;k3E0PDA�TE P��?KS_24�1G��_INFO 1+������10%  �OLGE011 y.��0056�� �5�G�*�k�}�`ߡ� �����ߺ������1���U�g�9��OFF�SET .�= q�l��0s�����������!�N�E�W����n�`����������� ��"O~��?{�
c2m?���UFR?AME  f5�����RTOL_AB�RT����ENB���GRP 1/��9�1Cz  A�:8l�8J\n������
�0U����MSK  �f5���	N�%���%KH/�2VCC�M��0��]"MR� 26T9 �e9�	��O�~�XC'�*�/�&X��� �5��A@�p��L. j8?d�7?I?v?Ч!q?�?5�A��l��?�?l�� B����1l��5�?Ob? ?OOcONO�OrO�O�O �O�O8O�O___M_  Oq_�_d���!�/�_ �/�/�/??'?o�O \oSo1_�o�o�?�?�o �?__�o"io{o=j U�y���-� ��	�B�U_f�x��� ��!�_���_�_�_o o'o��\�S�1��� ���o�oڟ�o_���"� i�{�=�j�U���y��� ��֯-���ɯ�	�B� U�f�x����=����� ͏ߏ���'��� \�S�1��ϤϷ�ɟ�� �_���"�i�{�=�j� Uߎ�y߲ߝ���-��� ���	�B�U�f�x�O/�ISIONTMOiU� $r%����d#7�K ��LT/ FR�:\��\DATA�\�� �� �MC��LOG�� �  UD1��E�X��' B@ ��O� �7/�m� �q���� ��  =	 1�- n6  -#��T�L�&,������=�����T����TRAIN�6������"8�+ (:���S.�Sa s��������'9KX&LE�XE��9�+�!1-�eR,MPHASE'  k%�#�R]!�SHIFTMEN�U 1:�+
 <a\�6//����� !/Z/1/C/�/g/y/�/ �/�/�/?�/�/D??�-?z?Q?	LIV�E/SNAPn3?vsfliv��?�^3�� SETU<�0�2menu�?�?�d?)O;OB��;����	(H'O�O\����� ��@�AV�B8`�`����H���A�B��C��G g��KSFME�0ة���� �MOڒ<��z��WA�ITDINEND���Q@WOK  !�X[]��w_S�_^YwTIM�����\GH_�]j_�[�_�Z�_x�Z�_\XRELE�`gU@T����AS_ACT�0
h�a\X�_�� =��b%�  OLGE12�5.	r0001<��bRDIS�0�o~APV_AXSRG`2>bJ<��O��Gp~4 _IR  � �᥀������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2��D�V�h�z�����ZA�BC31?bI�� 	,�=�2��ܬ¯������
��Y���MPCF_G 1@S}0A�������ҿ�������,�b�MP��A�bI  �@���8:��Q8|O��0��t��Ϙ�?�T��� ����D����k�-ߞ����ѿp��������� ��	�l�E��i�{�� ��R�\�n߀ߚ���� ��2���e�w���� ������.��d�= OZ�s�@��\� ����'9���� Tf�����& �/5/�\// �/B/T/f/x/�/�/F ��(?:?L?v>��u��(PBS{j�P_CY�LINDER 2�CS{ ��& ,(  *�?�=�#`�?O�?8OM �/ nO�O�N�?�O$O�O�O �O_RO3_E_W_�O{_ _�O�_�_�_�_*_o�of�R�2DSw�a �"�hoxl�s�/�o@�o�o��o�o�1�qA��o*yo�o`�o ��o}�	��? y&�uJ��Z���� m����?��׏�_��4�F����2SPHE_RE 2E�=�o_ ���_��͟����_L� '�9�i_]���⟓�z� ��������F�X�5� ��Y�@�R���֯��ſ|׿N�ZZ  �$��4