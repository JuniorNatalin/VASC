��   t��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���U�I_CONFIG�_T  d �9$NUM_MENUS  9�* NECTCRE�COVER>CCOLOR_CRR�:EXTSTAT���$TOP>_�IDXCMEM_�LIMIR$D�BGLVL�PO�PUP_MASK��zA  $DUMMY54��ODE�
5CFO�CA �6CPS�)C��g HA�N� � TIME�OU�PIPES�IZE � MW�IN�PANEM;AP�  � � �FAVB ?� 
w$HL�_DIQ�?� qELEM�Z�UR� l� S|s�$HMI��RO+\W AD�ONLY� �T�OUCH�PRO�OMMO#?$��ALAR< �F�ILVEW�	E�NB=%%fC �1"USER:)FC[TN:)WI�� I* _ED�l"V!�_TITL� ~1"COORDF<#/LOCK6%�$F%|�!b"EBFOR�? �"e&
�"�%�!�BA�!j ?�"B�G�%$PM�X�_PKT�"IHE�LP� MER�B�LNK$=ENAB��!? SIPMAN�UA�-4"="�B�EEY?$�=&q!E�Dy#�&UST�OM0 t �$} RT_SPI�D��4C�4*PA�G� ?^DEV�ICE�9SCREVuEF���7N��@$FLAG�@��&�1  h� 	$PWD_A�CCES� E �8��TC�!�%)$�LABE� 	$	Tz j4@q!�D��	L&USRV�I 1  < �`� �B��APRI�m� U1�@�TRIP�"m�$�$CLA?@ �����A��R��R��$'2 ~����R�	 �,��?���/Q�>P8R3T.Q��	���)P�  �?����
 ���A�_�_�_�_�_�_o �_*o<oNo`oro �oo�o�o�o�o�o �o&8J\n����(/SOFTP��0/GENLIN�K?curren�t=menupa�ge,935,1 �����!:�L� ^�p�����#���ʏ܏ � ����6�H�Z�l� ~�����1�Ɵ؟��� � ���D�V�h�z�������� TPTX����:�ٯ��� s Ƿ����$/softpa�rt/genli�nk?help=�/md/tp�q.dg��F�X�j�|�5�9&�#�pwd2�ɿ ۿ���4�#�5�G�Y� k�}�ϡϳ������� �ϊϜ�1�C�U�g�y�T��aT��AsVQR�� ($ �����`�����(����A�2QN�PS2S������D�^�
q�2QtQ��,RQ  ��ʡSV�������L�L�rY�S�2 1�E~>PR \ �}mPRE�G VED��6�H��wholemod�.htm\�sin�glm�doub~��trip��brows�� ��I�������3E Wi{�3�W�i�_dev.sr�l�4��	1�	t �� 	��o��]������(/�  �@@/R/d/v/�/�/�/0�/�/�/�& @</? #?�/G?Y?k?:6+�#/ /�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O��O�O#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCo Uogo5/�o�o�o�o�o �o 2D??hz I[��y?�?qo
� ��)�R�M�_�q��� �������ݏ��*� %�7�_W�Q������ ��ǟٟ����!�3� E�W�i�{�������ï �o���"�4�F�X�j� |������Ŀֿ���� ����ͯf�a�s� �Ϯϩϻ�������� �>�9�K�]߆߁ߓ� a��߭��������#� 5�G�Y�k�}���� �����������Z� l�~������������� ���� 2hz 1�C�)�����
 )RM_q� ��������/ 	/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?I��?�?�? �?�?O"O4OFOXOS�|O�O]OoO�O�O�J��$UI_TOPMENU 1�@�QR 
�XQ�1)*d?efault�?�=�	*levelw0 *HP 8_�& o__m_Rtp�io[23](?tpst[1�X�_��_�_BVX_�_!$
h�58e01.gi�fo(	menu15Bi9`da13Bjcb�Ajad4ikPoa�� �o�o�o $6�2 �o_q����Ht�prim=dap�age,1422,1����/�A� Le�w���������N���vclass,5ȏ���!�3�E�P�܌13L�������h��ʟQ��|53�@��*�<�N�Q��|8����������ѯP������+�=�O��9 PQ_��B]y�aw��oÿ�Vty�]�_�QOmf[0�_��	�c[164�W>�5�9�Xa�oٿ{�]h2 �ogm��}j�osgAk�� �cg�y�F�X�j�|ߎ� 寲����������� 0�B�T�f�x���ۍ2������������ �O�a�s�����&�8� p������� ۟�14�^p���%���sainedi����%�wintp�p0bt ����6Qr��� fo��//0/B/T/ f/x/�/ o�/�/�/�/ �/??,?>?c?�o�? �?�?�?�?�? �OO )O;OMO_O�?�O�O�O �O�O�O�O~O_%_7_ I_[_m_�O�_�_�_�_ �_�_z_o!o3oEoWo io{o
o�o�o�o�o�o �o�o/ASew ��������o�0������⯿]?o��s󽌏������u��d�f���&�4�@���B�h��ό�6��u7���0���� '�9��]�o������� ��F�ۯ����#�5�G�64�1C����� ����ɿԯ����#� 5�G�ֿk�}Ϗϡϳ� ����2�����1�C�U�����6\ߑߣߵ�0����4Ӝ74�� '�9�K�]������ �/z����������"� G�F���R�|������� ��������p?1CU gy�Vϯ��� �	�?Qcu ��(����/ /�;/M/_/q/�/�/ �/6/�/�/�/??%? �/I?[?m??�?�?2? �?�?�?�?O!O3O�? WOiO{O�O�O�Ol�~� �O��l�
_._@_R_ w_v_�_�__�_�_�_ ooo*o<oNo�o �o�o�o�o�o�oHO '9K]o�o�� ����|�#�5� G�Y�k�}������ŏ ׏������1�C�U� g�y��������ӟ� ��	���-�?�Q�c�u� �������ϯ��� �O�O;��O�_^op��� ������ʿܿ�\��� 7�6�H�Z�l�~ϐϢ� po�������!�3�E� ��i�{ߍߟ߱���R� ������/�A�S��� w�������`��� ��+�=�O���s��� ����������n� '9K]����� ���j�#5 GYk&����ϲ� ����//0/B/ �b/`/�/�/�/�/�/ �/�/?��??Q?c?u? �?�?��?�?�?�?O O�?;OMO_OqO�O�O �O6O�O�O�O__%_ �OI_[_m__�_�_2_ �_�_�_�_o!o3o�_ Woio{o�o�o�o@o�o �o�o/�oSe w����z�� �??*�<�N�`�r� ���������ޏ��� �&�K�J�\�*?���� ��ɟ۟�D�#�5� G�Y�k�}������ů ׯ������1�C�U� g�y��������ӿ� ��	Ϙ�-�?�Q�c�u� ��ϫϽ�������� ��)�;�M�_�q߃ߕ� $߹����������w��t*defau�lt�w�*level8ˏi�{���7� tpst�[1]����y��tpio[23������u��n��6�H��	menu7.gkifI�
h�13m�Bz�5��g��e�4��u6m�����% 7I��m��� �V��!3E�W�prim=�h�page,74,1\�������pclass,13�/(/:/L/^/��5d/�/�/�/�/�/���/?.?`@?R?d?gy18���?�?�?�?�?�/�6��?%O7OIO[OmOL���$UI_USERVIEW 1�q��qR 
��tON�O�OF�m�O__%_7_I_ �Om__�_�_�_X_�_ �_�_o!o�O.o@oRo �_�o�o�o�o�oxo�o /AS�ow� ���jo���b +�=�O�a�s������ ��͏ߏ����'�9��K��*zoom>^�ZOOM]�� ��ԟ���
���.� @�R�d�v���������Я���*ma�xres��MAXRES������\� n�������G�ȿڿ� ��ϳ�4�F�X�j�|� '��ϛϭ������� �0�B���f�xߊߜ� ��Q����������� '�=�K�߆���� ��q�����(�:�L� ��p���������c��� ����[�$6HZl �����{�  2D��Ucu ������
/� ./@/R/d/v//�/�/ �/�/�/��/??�/ N?`?r?�?�?9?�?�? �?�?OO�?8OJO\O nO�O#A