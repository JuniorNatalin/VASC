��   �P�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�RYRUN_T   � $'�ENB 4 NU�M_PORTA �ESU@$ST�ATE P TC�OL_��PMPM�CmGRP_MA�SKZE� OTI�ONNLOG_IgNFONiAVc�FLTR_EMP�TYd $PRO�D__ L �ESTOP_DSBLA�POW_RECO�VAOPR�SA�W_� G %�$INIT	RE�SUME_TYP�EN@&J_ � 4 $($FST_IDX��P_ICI |�MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI��.yMKR-�  $LIN�c   �_SIZc�x� k�. , $USE_FL4 �p�&i*SIMA��Q#QB6'SC�AN�AXS+IN�S*I��_COUN�rRO��_!_TMR_VA�g�h>�i) �'�` ��R��!�+W[AR�$}H�!�{#NPCH���$$CLASS ? ���01���5��5�6/ 05�5�����c"����\1l51071|p5��%VAG4���<�0TP�?���A5I2L;cK ��"��	A$��Y4d��Y3	A[2�)Y3�Y4-D *&H��&G\0pA�hF	~ChF�ChF�T�ChF�n@�fH̾C�hF�n@�fH�n@��&GAA4B�D!z08P�H`0Q�Fhz0i�H�l.S�Fyz0��H��z0��H�z0��H��z0�&G~SxV�~P�HU@�QxVa@U2vX9~P;vXA~PUPvXa~PxvX��S*xV�~P�vX�cxVe�~P�vX�@�vX��>cxV�~P�@xV�^c(E\0Phf=@K+fhC�chfH# ��5maL�chfQ# q,fhAP{fh��chf�# QPhf��chfaP�qPhf�@�fh�L# Eh�>s(E�@XPqHvP3Fx7ns`Hv�0�qHv�PsFx�w�sHv��sHv!`Y�Fx1p�&G�@$�q�v �s�v1�p�P��vV�p�P�vv�p�T��=AD��G&�M��X�U=AAP z&�^�*)�����&��~�)���q�&����&��B��&�ae=A���(eU=A�A�&����@(� ��P����P ���J.����P @����PP���` U��en���u �U���U������ �&�
n@�P(���DB���z0��?���������6W?05�V1 FOwLGE��U�U~e�MAKROq��SUCH�eh�B�IN���*�`��o { 2L; 74%|�SP��֯z���J�Z5Ʀ<�U
�  Ne�q��6Ʀeu>�  na%m�}1Ʀ4A���� v�Y�;2����1�"-��̠6����m� n��̠uu�  ter�̠UB�@-��%�����L?�ʁ�����PA ����X �01\0s2�tq* Z����t�����=��t ���� E����#�5�G�Y�k� }ߏߡ�����p6}1�������(tOq
_Pqu��Q��Rt��}1	��-�?� Q�c�u�����71���&Ū�!2t�� �����d�ss��k��p��n���o�tr
 ��8�J�\�n�����@������������&��Wds��k��p��n��o'�>Pb t�������
��$���� ASew����P�����)��� $6N/`/r/�/�/�/@�/�/�/�/?��(����=/O?a?s?�? �?�?�?�?�?�?O��!��O;OMO_OqO�O �O�O�O�O�O�O__l����d�C��DB?S_e_w_�_�_ �_�_�_�_�_oo����:P>_Woio {o�o�o�o�o�o�o�o (o+Sew� ���������+�&\
6Q )�� +T�7Joo������� ��ɏۏ����#�5���>_�q������� ��˟ݟ���%�7� :�D�k�}�������ů ׯ�����1�C�N� g�y���������ӿ� ��	��-�?�Q�\�u� �ϙϫϽ�������� �)�;�M�X�\߃ߕ� �߹���������%� 7�I�[�f����� ���������!�3�E� W�i�t���������� ����/ASe p�t������ +=Oas~ ������// '/9/K/]/o/�/��/ �/�/�/�/�/?#?5?�G?Y?k?}?�/2Pd�s2Pq2P!�1#
�1%�1'^��?�?�? OO+O=OOOaOsO�O*@�F��7"�?�O �O�O __$_6_H_Z_Pl_~_�_�O�L$�O �_�_�_oo1oCoUo�goyo�o�o�J�2  �_�_�o�o/A�Sew���oH� �l�O��
��.�@��R�d�v��������K.� &�1(��� ��/�A�S�e�w����������0�?���� ��/�A�S�e�w��� �������Eï���� !�3�E�W�i�{����� ��ÿ�/�����/� A�S�e�wωϛϭϿ���Ϝ6ds
 q���
��.� @�R�d�v߈ߚ߬߾���ߔ7�t��Ckqu��D��E��UF�G��H��I�Jt��5�G�Y�k�}�@����������2�tW ds��C�D��UE�F��G�H�I��"�;�M�_�q��� ������������1��UK��L�M��N�UO��P�Q��R,� DVhz����������p��K�L���M�N��O�P��Q�2K]o� ��������q
��S��T;3/E/W/ i/{/�/�/�/�/�/�/T�/�6�t$��S� !/:?L?^?p?�?�?�?@�?�?�?�? O?%��UU%1V��W%1X*? NO`OrO�O�O�O�O�OP�O�O_���t&��U��V%1W��<OU_ g_y_�_�_�_�_�_�_P�_	o_�t'��Y%1Z��[%1\E_^opo �o�o�o�o�o�o�o �oǃ(��Y��Z%1[��Loew�� �������$>4)ds2 U[� m��������Ǐُ�P���!���	4*F� _�q���������˟ݟ@���%�7�B�+N� g�y���������ӯ�@��	��-�?�B�,V� o���������ɿۿ�@���#�5�G�B�-^� wωϛϭϿ�������@��+�=�O�B�.f� ߑߣߵ���������@�!�3�E�W�b�/n� ������������@�)�;�M�_�b�0v� ��������������@1CUgb�1~� ������@'9K]ob�2� ������//@//A/S/e/w/b�3� �/�/�/�/�/??%?@7?I?[?m??b�4�/ �?�?�?�?�?	OO-O@?OQOcOuO�Ob�5�? �O�O�O�O�O_#_5_@G_Y_k_}_�_b�6�O �_�_�_�_oo+o=o@Ooaoso�o�ob�7�_ �o�o�o�o!3E@Wi{��b�8�o �����)�;�M�@_�q��������x9� ׏�����1�C�U�@g�y��������x:Ə ߟ���'�9�K�]�@o����������x;Ο �����/�A�S�e�@w����������x<֯ ���%�7�I�[�m�@ϑϣϵ��ϲx=޿ ��	��-�?�Q�c�u�@�ߙ߽߫��߲x>�� ���#�5�G�Y�k�}�@��������x?�� ��+�=�O�a�s���@�����������x@�� !3EWi{�@������xA�� );M_q��@������xB /1/C/U/g/y/�/�/@�/�/�/�/�/�xC/ '?9?K?]?o?�?�?�?@�?�?�?�?�?�xD? /OAOSOeOwO�O�O�O �O�O�O�O_�u_3_ E_W_i_{_�_�_�_�_ �_�_�_o�u_7oIo [omoo�o�o�o�o�o �o�oo3EWi {������� ��(A�S�e�w��� ������я����� +�6�O�a�s������� ��͟ߟ���'�2� K�]�o���������ɯ ۯ����#�5�@�Y� k�}�������ſ׿� ����1�C�N�g�y� �ϝϯ���������	� �-�?�J�c�u߇ߙ� �߽���������)� ;�M�X�q����� ��������%�7�I� [�f������������ ����!3EWb� {������� /ASep� ������// +/=/O/a/s/~�/�/ �/�/�/�/??'?9? K?]?o?z/�?�?�?�? �?�?�?O#O5OGOYO kO}O�?�O�O�O�O�O �O__1_C_U_g_y_ �_�O�_�_�_�_�_	o o-o?oQocouo�o�_ �o�o�o�o�o) ;M_q���o� �����%�7�I� [�m�������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ư߿���'�9� K�]�oρϓϥϷ�¿ �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q��������� `ds2t�&8J \n������ ���/"/4/F/X/j/ |/�/�/�/�/�/�/� ??0?B?T?f?x?�? �?�?�?�?�?�??O ,O>OPObOtO�O�O�O �O�O�O�O�?O(_:_ L_^_p_�_�_�_�_�_ �_�_ o_$o6oHoZo lo~o�o�o�o�o�o�o �oo2DVhz �������
� '@�R�d�v����� ����Џ����#� <�N�`�r��������� ̟ޟ���&�1�J� \�n���������ȯگ ����"�-�?�X�j� |�������Ŀֿ��� ��0�;�T�f�xϊ� �Ϯ����������� ,�>�I�b�t߆ߘߪ� ����������(�:� E�W�p������� ���� ��$�6�H�S� l�~������������� �� 2DVa�z �������
 .@R]o�� �����//*/ </N/`/k�/�/�/�/ �/�/�/??&?8?J? \?n?y/�?�?�?�?�? �?�?O"O4OFOXOjO u?�?�O�O�O�O�O�O __0_B_T_f_x_�O �_�_�_�_�_�_oo ,o>oPoboto�o�_�o �o�o�o�o(: L^p��o�o�� �� ��$�6�H�Z� l�~������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲߽������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p����� ���� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�
? ?.?@?R?d?v?�?�? �?�?�?�?�/�/O*O <ONO`OrO�O�O�O�O �O�O�O�?_&_8_J_ \_n_�_�_�_�_�_�_ �_�_	_"o4oFoXojo |o�o�o�o�o�o�o�o oo0BTfx� ������� ,�>�P�b�t������� ��Ώ�����!�:� L�^�p���������ʟ ܟ� ���/�H�Z� l�~�������Ưد� ��� �+�D�V�h�z� ������¿Կ���
� �.�9�R�d�vψϚ� �Ͼ���������*� 5�G�`�r߄ߖߨߺ� ��������&�8�C� \�n��������� �����"�4�F�Q�j� |��������������� 0BM�_�x� ������ ,>P[t��� ����//(/:/ L/^/i�/�/�/�/�/ �/�/ ??$?6?H?Z? e/w/�?�?�?�?�?�? �?O O2ODOVOhOs<�* �ds
��r
 t tO�O�O�O�O�O__@)_;_M___q_u6~? �_�_�_�_�_�_oo /oAoSoeowor?�o�o �o�o�o�o+= Oas��o��� ����'�9�K�]� o��������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϲ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ���'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/��/? ?1?C?U?g?y?�?�? �?�?�?�?�/	OO-O ?OQOcOuO�O�O�O�O �O�O�O�?_)_;_M_ __q_�_�_�_�_�_�_ �_�Oo%o7oIo[omo o�o�o�o�o�o�o�o o!3EWi{� ������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ��� �9�K�]� o���������ɯۯ� ���#�.�G�Y�k�}� ������ſ׿���� �*�C�U�g�yϋϝ� ����������	��-� 8�Q�c�u߇ߙ߽߫� ��������)�;�F� _�q��������� ����%�7�B�[�m� ��������������� !3EP�i{� ������ /AS^w��� ����//+/=/ O/Zs/�/�/�/�/�/ �/�/??'?9?K?]? h/�?�?�?�?�?�?�? �?O#O5OGOYOkOv? �O�O�O�O�O�O�O_ _1_C_U_g_rO�_�_ �_�_�_�_�_	oo-o ?oQocouo�_�o�o�o �o�o�o);M _q��o���� ���%�7�I�[�m� ������Ǐُ��� �!�3�E�W�i�{��� ����ß՟����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϰ������� ���#�5�G�Y�k�}� �ߡ߳߾�������� �1�C�U�g�y��� ���������	��-� ?�Q�c�u��������� ������);M _q������� �%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/��/?? /?A?S?e?w?�?�?�? �?�?�?�/OO+O=O OOaOsO�O�O�O�O�O �O�?__'_9_K_]_ o_�_�_�_�_�_�_�_ �Oo#o5oGoYoko}o �o�o�o�o�o�o�oo 1CUgy�� ������-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ����7�I�[�m� �������ǯٯ��� ��3�E�W�i�{��� ����ÿտ����� (�A�S�e�wωϛϭ� ����������+�