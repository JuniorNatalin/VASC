��   �P�A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�RYRUN_T   � $'�ENB 4 NU�M_PORTA �ESU@$ST�ATE P TC�OL_��PMPM�CmGRP_MA�SKZE� OTI�ONNLOG_IgNFONiAVc�FLTR_EMP�TYd $PRO�D__ L �ESTOP_DSBLA�POW_RECO�VAOPR�SA�W_� G %�$INIT	RE�SUME_TYP�EN,&J_ � 4 $($FST_IDX��P_ICI��MIX_BG-yA
_NAMc �MODc_US�d�IFY_TI� �xMKR�-  $L{INc   �o_SIZc@x�� k. , $USE_FL�4 ��&i*SIAMA�Q#QB6'oSCAN�AXS+�INS*I��_COUNrRO��_!_TMR_VA�g�h>�i ) �'` ��R��!n�+WAR�$}iH�!{#NPCH���$$CLAS�S  ���401��5��5�6/ �055���c*����i81071>��%VAG�?�<�0TP�?���A5I2L;c ���"��	A$���m4d��m3	Ao2)fm3�m4-D &H��&Gp0pAhFI	~ChF�ChFÞC*hF�n@�fH̾ChFU�n@�fH�n@�&GQAA4B�D!z08�H�`0Q�Fhz0i�HlT.S�Fyz0��H�z0U��H�z0��H�z0M�&G~SxV~PHU@�QxVa@2�vX9~P;vXA~PP*vXa~PxvX��SxV��~P�vX�cxV��~P�vX�@�vX�D>cxV�~P�@xV�^c�(Ep0Phf=@%+fhC�chfH# �5RmaL�chfQ# qfh�AP{fh��chf��# QPhf��chfaPXqPhf�@�fh�# &Eh�>s(E�@Pq,HvP3Fx7nsHv��0�qHv�PsFxwĞsHv��sHv!`�,Fx1p�&G�@�q�v �s�v1�p�P�vQV�p�P�vv�p���*=AD��G&�M���U,=AAP z&�^�)�����&��~�)��qU�&����&����!�&�ae=A���eU=A�A�&����@(� ��P����P ���J.����P@����PP���` U��	en���u �U��U�Ԑ���� �&�
�n@�P(���DB���z0��?�������l�6W?05V1� FOL�GE��U�U � 0h�MAKR}Oa�SUCH�e�h�BIN���sD�o { 2L;� 4%|�SP蟦ׯ���J{���Ʀ�U
�  </�t�̠eu>�  hI=eq%�}1Ʀ4A���5-��Y�;2����="k���6���\�<uu�  amu���UB����"�����L=p1�������PXA ��%�X �01�p0s* q����� ��!��_&��`t����t��F� ��'�9�K�]�o߁��ߥ���m9}1����Bqu) H�ҷIqs��Zr��\�ttq�иttt }1�'�9�K�]�o�� ��������UA�0� 2L9 ������dss
�^q	�_tr
 t��*�<� N�`�r����������������@��dsu	�_�,>Pb t������� ��?o6*<N` r������� /0A*/</N/`/r/ �/�/�/�/�/�/�/? /&?8?J?\?n?�?�? �?�?�?�?�?�?O? 4OFOXOjO|O�O�O�O �O�O�O�O_O)OB_ T_f_x_�_�_�_�_�_ �_�_oo%_>oPobo to�o�o�o�o�o�o�o (3oL^p� ������ �� $�/AZ�l�~����� ��Ə؏���� �2� =�V�h�z������� ԟ���
��.�@�K� d�v���������Я� ����*�<�G�Y�r� ��������̿޿�� �&�8�J�U�nπϒ� �϶����������"� 4�F�X�c�|ߎߠ߲� ����������0�B� T�_�qߊ������� ������,�>�P�b� m�������������� (:L^p{� ������  $6HZlw�� �����/ /2/ D/V/h/z/��/�/�/ �/�/�/
??.?@?R? d?v?�?�/�?�?�?�? �?OO*O<ONO`OrO �O�?�?�O�O�O�O_ _&_8_J_\_n_�_�_ �O�_�_�_�_�_o"o 4oFoXojo|o�o�o�_ �o�o�o�o0B Tfx���o�o� ����,�>�P�b� t��������Ώ��� ��(�:�L�^�p��� ������Ïܟ� �� $�6�H�Z�l�~����� ����џ���� �2� D�V�h�z�������¿ ͯ���
��.�@�R� d�vψϚϬϾ���۴�* ds
� q����t���"�4�F�X�j߀|ߎߠ߲�����ڱz����Cqu��UD��E��F��G��UH��I��J��K��L��?�Q�c�u��ﰫ������ =�� �ds��C��D��E���F��G��H��I
��J��K��-�F�X� j�|����������������!��M��N��O��P6�/ASew�����������"��6H Zl~����������#ds2  &+/=/O/a/s/�/�/@�/�/�/�/�/��	��$//?A?S?e?w?�? �?�?�?�?�?�?O8%?7OIO[OmOO�O �O�O�O�O�O�O_8&&O?_Q_c_u_�_�_ �_�_�_�_�_oo8'._GoYoko}o�o�o �o�o�o�o�o8(6oOas��� ������'�8)>W�i�{������� ÏՏ�����/�8*F�_�q��������� ˟ݟ���%�7�8+N�g�y��������� ӯ���	��-�?�8,V�o���������ɿ ۿ����#�5�G�8-^�wωϛϭϿ��� ������+�=�O�8.f�ߑߣߵ����� �����!�3�E�W�b�/n߇�������� ����)�;�M�_�b�0v������������ ��1CUgb�1~������� '9K]ob�2������� ////A/S/e/w/�3��/�/�/�/�/? ?%?7?I?[?m??�4�/�?�?�?�?�?	O O-O?OQOcOuO�O�5�?�O�O�O�O�O_ #_5_G_Y_k_}_�_�6�O�_�_�_�_oo +o=oOoaoso�o�o�7�_�o�o�o�o! 3EWi{���8�o�����)� ;�M�_�q��������9�׏�����1� C�U�g�y��������:Əߟ���'�9� K�]�o����������;Ο�����/�A� S�e�w����������<֯���%�7�I� [�m�ϑϣϵ��ς=޿��	��-�?�Q� c�u߇ߙ߽߫��߂>�����#�5�G�Y� k�}��������?����+�=�O�a� s��������������@��!3EWi {�������A��);M_q ��������(B/1/C/U/g/y/ �/�/�/�/�/�/�/(C/'?9?K?]?o?�? �?�?�?�?�?�?�?(D?/OAOSOeOwO�O �O�O�O�O�O�O_% _3_E_W_i_{_�_�_ �_�_�_�_�_o�_ 7oIo[omoo�o�o�o �o�o�o�oo3E Wi{����� ����(A�S�e� w���������я��� ��+�6�O�a�s��� ������͟ߟ��� '�2�K�]�o������� ��ɯۯ����#�5� @�Y�k�}�������ſ ׿�����1�C�N� g�yϋϝϯ������� ��	��-�?�J�c�u� �ߙ߽߫�������� �)�;�M�X�q��� �����������%� 7�I�[�f�������� ��������!3E Wb�{����� ��/ASe p������� //+/=/O/a/s/~ �/�/�/�/�/�/?? '?9?K?]?o?z/�?�? �?�?�?�?�?O#O5O GOYOkO}O�?�O�O�O �O�O�O__1_C_U_ g_y_�_�O�_�_�_�_ �_	oo-o?oQocouo �o�_�o�o�o�o�o );M_q�� �o������%� 7�I�[�m������� Ǐُ����!�3�E� W�i�{�������ß՟ �����/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ư߿��� '�9�K�]�oρϓϥ� ��¿�������#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u��������������*� _ds
�[qu���q�����qss�����tr t��6 q �t��C Ugy�����j��@��`��J �L K Mqu�qs)Ar�skq)� �t!'�tt1K]o���������A��akds���,�rK8tB,  u(�H""I Z  \9J/\/n/�/�/�/ �/�/�/�/��9��? )?;?M?_?q?�?�?�? �?�?�?�?��O%O7O IO[OmOO�O�O�O�O �O�O�OO!_3_E_W_ i_{_�_�_�_�_�_�_ �_o_/oAoSoeowo �o�o�o�o�o�o�o o+=Oas�� �������  9�K�]�o��������� ɏۏ����#�.�G� Y�k�}�������şן �����*�C�U�g� y���������ӯ��� 	��-�8�Q�c�u��� ������Ͽ���� )�;�F�_�qσϕϧ� ����������%�7� B�[�m�ߑߣߵ��� �������!�3�E�P� i�{���������� ����/�A�S�^�w� �������������� +=OZ�s�� �����' 9K]h���� ����/#/5/G/ Y/k/v�/�/�/�/�/ �/�/??1?C?U?g? r/�?�?�?�?�?�?�? 	OO-O?OQOcOuO�? �O�O�O�O�O�O__ )_;_M___q_�_�O�_ �_�_�_�_oo%o7o Io[omoo�_�o�o�o �o�o�o!3EW i{��o���� ���/�A�S�e�w� �������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}���������׿ �����1�C�U�g� yϋϝϯϺ������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������� �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�??'? 9?K?]?o?�?�?�?�? �?�?�?�/O#O5OGO YOkO}O�O�O�O�O�O �O�OO_1_C_U_g_ y_�_�_�_�_�_�_�_ _o-o?oQocouo�o �o�o�o�o�o�oo );M_q��� ������7� I�[�m��������Ǐ ُ�����3�E�W� i�{�������ß՟� ����(�A�S�e�w� ��������ѯ���� �+�6�O�a�s����� ����Ϳ߿���'� 2�K�]�oρϓϥϷ� ���������#�5�@� Y�k�}ߏߡ߳����� ������1�C�N�g� y������������ 	��-�?�J�c�u��� ������������ );MX�q��� ����%7 I[f���� ���/!/3/E/W/ b{/�/�/�/�/�/�/ �/??/?A?S?e?p/ �?�?�?�?�?�?�?O O+O=OOOaOsO~?�O �O�O�O�O�O__'_ 9_K_]_o_zO�_�_�_ �_�_�_�_o#o5oGo Yoko}o�_�o�o�o�o �o�o1CUg y��o����� 	��-�?�Q�c�u��� �����Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϸ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y�������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�??%?7? I?[?m??�?�?�?�? �?�?�/O!O3OEOWO iO{O�O�O�O�O�O�O �?__/_A_S_e_w_ �_�_�_�_�_�_�_ _ o+o=oOoaoso�o�o �o�o�o�o�oo' 9K]o���� ����
#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��&�?�Q�c�u��� ������ϯ���� "�;�M�_�q������� ��˿ݿ���%�0� I�[�m�ϑϣϵ��� �������!�3�>�W� i�{ߍߟ߱������� ����/�:�S�e�w� ������������ �+�=�H�a�s����� ����������' 9KV�o���� ����#5G Rk}����� ��//1/C/U/` y/�/�/�/�/�/�/�/ 	??-???Q?c?n/�? �?�?�?�?�?�?OO )O;OMO_Oj?�O�O�O �O�O�O�O__%_7_ I_[_m_xO�_�_�_�_ �_�_�_o!o3oEoWo io{o�_�o�o�o�o�o �o/ASew �o������� �+�=�O�a�s���� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫ϶��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew �������� +=Oas�� �����//'/ 9/K/]/o/�/�/�/�/ �/�/��/?#?5?G? Y?k?}?�?�?�?�?�? �/�?OO1OCOUOgO yO�O�O�O�O�O�O�? 	__-_?_Q_c_u_�_ �_�_�_�_�_�_�Oo )o;oMo_oqo�o�o�o �o�o�o�o�_%7 I[m���� ���!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯��� � 9�K�]�o��������� ɿۿ����#�.�G� Y�k�}Ϗϡϳ����� ������1�