A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �UI_CONFIG_T  d 9$NUM_MENUS  $NUM_CONNECT  $RECOVERMENU  $COLOR_CRT  $NUM_EXTSTAT   $TOPMENU_IDX  $MEM_LIMIT  $DBGLVL  $POPUP_MASK  $EXTSTATUS   $DUMMY54  $MODE   $DUMMY55  $FOCUS   $DUMMY56  $PS_CONFIG_C   $CONFIG_CHAN   $TIMEOUT  $PIPESIZE  $MWIN_LIMIT  $PANEMAP   $MENU_FAVS ?� 
$HLPMEN_DICT ? $HLPMEN_ELEM   $HLPMEN_URL ?� $DSPMEN_MASK  $HMI_MASK  $ROTIMEOUT   $READONLY   $TOUCH_MASK  $PROG_COMMON ?$ $ALARM_MASK  $FILVEW_MASK  $PS_ENB_MENU   $ENB_MENUFAV  $ENB_USERFAV  $ENB_FCTNFAV  $ENB_WIDE   $ICON_EDIT   $FCTN_TITLE $ENB_COORDFV  $LOCKMENUFAV  $LOCKUSERFAV  $ENB_WEBFORM  $COORD_FAVS   
$LOCKCOORDFV  $BACKCOLOR  $LOCKBGCOLOR  $PMN_MAX_PKT  $IHELP_TIMER  $BLNK_TIMER  $BLNK_ENABLE  $SIPMANUAL  $BLNK_ALARM  $TOUCH_BEEP  $ENB_TOPMENU  $ENB_ICONEDT   �UI_CUSTOM_T  t $START_SPID  $START_SCID  $CONFIG_PAGE ? $DEVICE_PAGE ? $SCREEN_DEF   �$CONFIG_PANE   @$FLAGS   @a��UI_TOPMENU_T  h 	$PWD_ACCESS  $DUMMY8  $PS_DUMMY   $DUMMY  $TITLE )$LABEL 	$TEXT ? 	$ICON ? 	$URL ?� 	,�UI_USRVIEW_T  < $MENU $CONFIG $FOCUS $PRIM m$DUAL m$TRIPLE m�$$CLASS  ������   R    R�$UI_CONFIG  ~���R	 ,           �  �       �                       , �                                 
 ���                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  �(/SOFTPART/GENLINK?current=menupage,935,1                                                                                          ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                    TPTX      TPTX      �          �          �             s �        ��$/softpart/genlink?help=/md/tpmenu.dg                                                                                              �&/softpart/genlink?help=/md/tpmenpwd.dg                                                                                            ��                                                                                                                                  ��                                                                                                                                  ��                                                                                                                                   ��                              ($�                                      $�                                      $�                                            �                                                    �                              
                                	     ���                                     �$UI_CUSTOM 1������R \  }     RESERVED              RESERVED              wholemod.htm          singlmod.htm          doublmod.htm          triplmod.htm          browsmod.htm          �                      RESERVED              RESERVED              RESERVED              �                      �                      �                      �                      �                        RESERVED              RESERVED              wholedev.stm          singldev.stm          doubdev1.stm          	tdev1.stm             browsdev.stm          �                      RESERVED              RESERVED              RESERVED              �                      �                      �                      �                      �                       � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ @ ���������������������������������������������������������������� @ ����������������������������������������������������������������  }     �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                        �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                       � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ @ ���������������������������������������������������������������� @ ����������������������������������������������������������������  }     �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                        �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                       � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ @ ���������������������������������������������������������������� @ ����������������������������������������������������������������  }     �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                        �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                       � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ @ ���������������������������������������������������������������� @ ����������������������������������������������������������������  }     �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                        �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                       � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ @ ���������������������������������������������������������������� @ �����������������������������������������������������������������$UI_TOPMENU 1������R 
X���    )*default                                  	*level0 *  	                                       *default                             tpio[23]          tpst[1]           *default          *default                              	                                       
h58e01.gif                           	menu5.gif         
menu13.gif        	menu1.gif         	menu4.gif                             	 ��                                                                                                                                   �                                                                                                                                   �prim=menupage,1422,1                                                                                                              �                                                                                                                                   �prim=menuclass,5                                                                                                                  �prim=menuclass,13                                                                                                                 �prim=menupage,153,1                                                                                                               �prim=menupage,18,1                                                                                                                �                                                                                                                                   �����)*default                                  	*level1    	 *default                                                tpty[1]           tpio[23]          tpmf[0]           *default          	tptc[164]         	tptc[159]          	 	menu4.gif                                               	menu2.gif         	menu5.gif         	menu3.gif         	menu1.gif         
menu11.gif        
menu11.gif         	 ��prim=menupage,18,1                                                                                                                �                                                                                                                                   �                                                                                                                                   �prim=menuclass,2                                                                                                                  �prim=menuclass,5                                                                                                                  �prim=menuclass,3                                                                                                                  �prim=menupage,151,1                                                                                                               �prim=mainedit                                                                                                                     �prim=wintpe,1                                                                                                                     ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �����)*default                                  	*level2    	 *default                                                tpsy[1]                                                 tpio[23]          tpsu[1]           *default           	 	menu4.gif                                               
menu15.gif                                              	menu5.gif         	menu6.gif         	menu7.gif          	 ��prim=menupage,18,1                                                                                                                �                                                                                                                                   �                                                                                                                                   �prim=menuclass,15                                                                                                                 �                                                                                                                                   �                                                                                                                                   �prim=menuclass,5                                                                                                                  �prim=menuclass,6                                                                                                                  �prim=menupage,74,1                                                                                                                ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   ������)                                           	            	                                                                                                                                                                             	                                                                                                                                                                             	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �                                                                                                                                    �����)*default                                  	*level8    	                                                          *default          tpst[1]           tpsy[1]           tpio[23]          *default          tpsu[1]            	                                                          	menu7.gif         
menu13.gif        
menu15.gif        	menu5.gif         	menu4.gif         	menu6.gif          	 ��                                                                                                                                   �                                                                                                                                   �                                                                                                                                   �prim=menupage,74,1                                                                                                                �prim=menuclass,13                                                                                                                 �prim=menuclass,15                                                                                                                 �prim=menuclass,5                                                                                                                  �prim=menupage,18,1                                                                                                                �prim=menuclass,6                                                                                                                  �$UI_USERVIEW 1������R 
��                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              *zoom                 ZOOM                  �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              *maxres               MAXRES                �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              �                      �                      �                      m�                                                                                                              m�                                                                                                              m�                                                                                                              