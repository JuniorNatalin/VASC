A��*SYSTEM*   V8.2306       4/24/2014 A   *SYSTEM*  �DRYRUN_T   � $DRYRUN_ENB  $NUM_PORT  $NUM_SUB  $STATE  $TCOL_SYSPT  $PMC_SYSPT  $GRP_MASK  $STEP_MOTION  $LOG_INFO  $TCOL_SAVE  $FLTR_EMPTY  $PROD_START  $ESTOP_DSBL  $POW_RECOV  $OPR_DSBL  $SAW_PROG %$INIT_PROG %$RESUME_TYPE  �DRYRUN_PORT_  4 $TYPE  $FST_IDX  $LST_IDX  $STATIC_PORT  ��MIX_BG_T  4 $PROG_NAME %$MODE  $STATUS  $MODIFY_TIME  �MIX_MKR_T   $LINE   $LINE_SIZE  �MIX_LOGIC_T , $USE_FLG  $USE_MKR  $USE_TCOL  $USE_TCOLSIM  $NUM_FLG  $NUM_MKR  $NUM_BG  $NUM_SCAN  $MAXNUM_SCAN  $MINNUM_SCAN  $ITEM_COUNT  $PROC_TIME  $MAX_TMR_VAL  $TCOL_LINE $TCOL_ENB  $TCOL_SIM  $TCOL_STAT  $SAVE_IDX  $SAVE_LINE $TCOL_WARN  $BG_HITEM  $INST_CHK  �$$CLASS  ������   5    5�$DRYRUN  ������5�      c                        ����                   %VAGSAW                                %VAGTPINI                                 �$DRYRUN_PORT 2������5� c    "      $             d                   )     �                                             	  	                    �  �         �  �         �  �         �  �         �  �                    !  8         c  c         h  i         l  l         y  �         �  �         �  �         �  �                      	                      2         9  ;         A  P         a  x         �  �         �  �         �  �         �  �         �  �         �  �         �  �         �  �           !         )  +         C  C         H  I         L  L         Q  q         y  {         �  �         �  �         �  �         �  �         �  �         �  �         �  �         	  	         !  3         7  7         I  I         a  s         w  w         �  �         �  �         �  �                                 1  A         V  a         v  �       )   D   G       )   M   P       )   y   z       )             )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )   �   �       )           )  !  !       )  2  2       )  J  J       )  A  A       )  P  P       )  `  c       )  e  e       )  u  x       )  z  z       )  �  �       )  
  9       )  �  �       )  �  �                                                                                                    �$DRYRUN_SUB ?������5�  FOLGE         UP            MAKRO      ) SUCHL         BIN1         x�$MIX_BG 2������5�  4%MAKROSP1                                    J� �%MAKROSP2                                    J� �%MAKROSP3                                    ����%MAKROSP4                                    ����%MAKROSP5                                    ����%MAKROSP6                                    ����%MAKROSP7                                    ����%MAKROSP8                                    J� ��$MIX_LOGIC ������5�                  �              X   ����  s2tq* q*  q* !q* #q* %q* 'q* )t* 't* $q* %t                                                                                                                                                                                                                     ����  * adss
�q�r)8tq
BqBqu) Hqu) Iqs) Zr) \ttq) �ttt�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   9          �$MIX_MKR 2������5 �  * dss
[q
]q
^q
_q
`tr
 tr
 t                                                                                                                                                                                                                       &  * dsu
[qu
]qu
^qu
_qu
`ttt`tt                                                                                                                                                                                                                        $  * dss
^q
_tr
 t
_qu
`tr
 tr
 t                                                                                                                                                                                                                         dss
Wqu
Xqu
]q
^q
_qu
`tr
 t                                                                                                                                                                                                                        * dss
[q
^q
_tr
 t
_q
`tr
 t                                                                                                                                                                                                                         * dss
]q
]q
^q
_q
`tr
 t                                                                                                                                                                                                                             &  * dss
]q
^q
_q
`tr
 t                                                                                                                                                                                                                                  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              * 
ds
 +q
 -t                                                                                                                                                                                                                                                     * dsu
 Aq
 Bt                                                                                                                                                                                                                                                    * ds
 Aqu
 Bt                                                                                                                                                                                                                                                    * ds* !q* #q* %q* )t                                                                                                                                                                                                                                           * dsu
 ?q
 @t                                                                                                                                                                                                                                                    * ds
 ?qu
 @t                                                                                                                                                                                                                                                    * dsu
 =q
 >t                                                                                                                                                                                                                                                    * ds
 =qu
 >r
 t                                                                                                                                                                                                                                               * dsu
 ;q
 <t                                                                                                                                                                                                                                                    * ds
 ;qu
 <t                                                                                                                                                                                                                                                    * dsu
 9q
 :t                                                                                                                                                                                                                                                    * ds
 9qu
 :t                                                                                                                                                                                                                                                    * ds
 )q
 /t                                                                                                                                                                                                                                                     * ds*  q* "t                                                                                                                                                                                                                                                     * ds* q* !t                                                                                                                                                                                                                                                     * ds* (q* *t                                                                                                                                                                                                                                                     * ds* 'q* )t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       * ds
 q
 t
t                                                                                                                                                                                                                                                * ds
Cqu
Dq
Equ
Ft                                                                                                                                                                                                                                         *  dsu
Cq
Dqu
Eq
Ft                                                                                                                                                                                                                                         * !ds
Gqu
Hq
Iqu
Jtt                                                                                                                                                                                                                                        * "dsu
Gq
Jqu
Iq
Jt                                                                                                                                                                                                                                         * #dsu
Kq
Lt                                                                                                                                                                                                                                                    * $ds
Kqu
Lt                                                                                                                                                                                                                                                    * %ds
Mqu
Nt
Mqu
Nt                                                                                                                                                                                                                                         * &dsu
Mq
Ntu
Mq
Nt                                                                                                                                                                                                                                         * 'dsu
Oq
Pru
Qq
Rtt                                                                                                                                                                                                                                        * (ds
Oqu
Pq
Qqu
Rtt                                                                                                                                                                                                                                        * )dsu
Sq
Ttu
Uq
Vt                                                                                                                                                                                                                                         * *ds
Squ
Tt
Uqu
Vt                                                                                                                                                                                                                                         * +dsu
Uq
Vt                                                                                                                                                                                                                                                    * ,ds
Uqu
Vt                                                                                                                                                                                                                                                    * -ds2 t                                                                                                                                                                                                                                                          	  * .ds2 t                                                                                                                                                                                                                                                          	  * /ds2 t                                                                                                                                                                                                                                                          	  * 0ds2 t                                                                                                                                                                                                                                                          	  * 1ds2 t                                                                                                                                                                                                                                                          	  * 2ds2 t                                                                                                                                                                                                                                                          	  * 3ds2 t                                                                                                                                                                                                                                                          	  * 4ds2 t                                                                                                                                                                                                                                                          	  * 5ds2 t                                                                                                                                                                                                                                                          	  * 6ds2 t                                                                                                                                                                                                                                                          	  * 7ds2 t                                                                                                                                                                                                                                                          	  * 8ds2 t                                                                                                                                                                                                                                                          	  * 9ds2 t                                                                                                                                                                                                                                                          	  * :ds2 t                                                                                                                                                                                                                                                          	  * ;ds2 t                                                                                                                                                                                                                                                          	  * <ds2 t                                                                                                                                                                                                                                                          	  * =ds2 t                                                                                                                                                                                                                                                          	  * >ds2 t                                                                                                                                                                                                                                                          	  * ?ds2 t                                                                                                                                                                                                                                                          	  * @ds2 t                                                                                                                                                                                                                                                          	  * Ads2 t                                                                                                                                                                                                                                                          	  * Bds2 t                                                                                                                                                                                                                                                          	  * Cds2 t                                                                                                                                                                                                                                                          	  * Dds2 t                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              * _ds
�qu
�q
�q
�qssu
�q
�tr�tqu
qu
q�t                                                                                                                                                                                                   @  * `ds
Jqu
Lqu
Kq
Mqu�qs)Arskq) �trsq) �ttt                                                                                                                                                                                                  A  * adss
�q�r)8tq
BqBqu) Hqu) Iqs) Zr) \tt                                                                                                                                                                                                          9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          