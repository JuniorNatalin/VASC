��   v��A��*SYST�EM*��V8.2�306 4/2�
 014 A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<�$1_8kW���FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\9 ^75z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D��VCAX_�w A.  @ 5vFX0OR�@E ?NUM_SE238�_TO0Q�#RE_:� 2cTW�+V>1 , $� �ME�vUPgDAT�wAXy_2 	T+VS5Q' 8<P��PnP;0k L\�R�PA�kQ�Q��+VM5Q  �$ISRTd 5+VG5Q { v��R2 
v�S2�T kR9�P 	��$U1SS  O����a����w�$' 1 �e� } �� 	 ����o�o�o�f�~����X��.u��5��� ����o�oA,s���p}���m ����
� �� ��F"���t�+w�a��}���� �{���:F�ʙ �Z ~Ь� ���|�+�=�d�a���p�� i7� uZ� ���wBB ���`B !��f�Xr��q(� ��fp�c~� ����o�7@�6_ `L�����% ����d�1�C�U����=L��`���?�����@���͟ߟ ���'�9�K�]�o������� �e��̧8��쯄d  2 �� /�A�S�e�w�����������<������ 1�C�U�g�yϋϝϯ� ���`�a�o������ *�<�#�`�K߄�oߨ� ��c��ߡ����&�[� 5�G�n�k�}����� ��������"���P� b�t������������� ��(:��^p ������Eϯ� �6HZl~� ����˿�/ / 2/D/V/h/z/�/�/�/ �/�/���/��/.?? R?9?v?a?�?�?�?�? ���?�?OO<O'O�? ]OoO�O�O�O�O3O�O �O_�O_J_=�k_}_ �_�_�_�_�_�_�_o o1oCoUo|o�o�o �o�o�o�goio�o- #Tfx���� �����,�>�P� b�t���������Ώ�� ��/�(��L�7�p� W������ʟ����? �՟6�!�Z�l��O{� ������ïկQ���� 2�D�/�h�[_������ ��ѿ�����+�=� O�a�s�5�ϬϾ��� ����G���'�K�A r߄ߖߨߺ������� ���m�J�\�n�� ����������������$FMS_G�RP 1^� >��J�|�H`k�G�SJ+4��H�MH�E9�J�2@�*Bu��C$26w���>��4��=�J�B�  ������IXB�������B#���±_�Bh���J���� N$ �Q��Q	Y�6LS1MN��:K�5f�@4���?����O�a�XJL��������\�*� �]  �} 	XJFE� ��� ��M.:S�M.;nM.<�N�6�N�v��N��N�Pg�O��O+1k�R�XS�g�s(s4s}V��Q�XJEJY�,�Y
-��Z�4��1���8��7.�3jp��3r��3����-H�-G���-F� ;޶��`�����-6���.�� ��-	�-(]���-��5�5�y�����������e����������������G���5�-P��-H��Hc�������n�� Q��*_���
�K �K ��������k��7 @�� ��U �f| ��d �ֶ ���� ��� ���@ �@  ��\U �tO ���f �� 0�u � ��3�� � l ��� 2�Hc"��	��y#��x-�u�������
������̰���]���f?������]J���>��4�� ��� �ǛS ��������M�!��M#�M�e�W���W����W��H�}���Jh���H�����W����T٥����_�X���X��G3�����q����c"���>C�"C���C�a7���7��7��� ����Dq���D�`�."��7��8D������7K_�7LI�0��1��7�� �'�c"  
�<d�4U��<�9�	��4�1T�4	��l4�F4��W�_�6  U(�B�A4��5z_��
������8
�	��4��*j�14���L@U��J4�~S@��NA������3�  |4�Y4��A3ᾪ@D����@�_�AgD3�n@@������KA�4�A\OCP  �4��4�UP�e4��,�4��h_��D�0��dFE�0�4o��.��kC�@��@z@����8,�D����_��[DNA*Q_��L@�,�vQ�(
�C�  +C�_��@��BXk#�_���3,4��oa�co7o�1)`�N�Aio{o�oT�4�%4�0�h;�hAh��c4�a�A54��Q�i�b8��{�;��8O��*�
��"�����s�M>j:I�?��	?��7�?��ӿ�m~����?e"�����ſ�������ʿ���?����(��7?��?���?��?�<��?�'5cs{�>�]?G�?m?<��?��5?� ������?���?�
`?����?��?_��?~��R�T�����n���*���þ��"���s�ɿ.̥��'��T ��]ž͝����!e� �K���_پ�Cξ��'������h�'
e�b�<�}?6�?�6�=?6ã?�7���Å>��B���rɿ��Z���p�?8�+�?9^6���?9]\?9�Y�+�"?9\m�<���G�+��b�P`��������� ����8_���?��Hy��8b���#z�����3C�ã������Ùb��߿â��è����������Or�q?���?��a?���?�3����>�����s��������7�?���?������?���Ӏ7?�u?����T,�?���	,($UP'004�o� ��4� �X�?�Q���u����� ���ϟ���a4����vA`�G�Y���}�.������7��毡�ߠ ��ȩ�Q��A���M�w� ^�������������ܹ23��'��K��o� Zϓϥϐ��ϴ����� ���5� �2�k�Vߏ� v߳ߞ�������� �+�=�gY�k�}�� �߳���T�������� 1�C�U�g�&������� ��������	��-? Qc"����| ���);M_ ����x�� /�%/7/I/[/// �/�/�/t/�/�/�/�/ !?3?E?W??{?�?�? �\a@p?�?�?�?d?O /OAOSOOwO�O�O�O lO�O�O�O�O_+_=_ O__s_�_�_�_h_�_��_�_�[��1234?567890o'e 	�oIo9omo]oyo�o �o�o�o�o�o�o! -5G{k��� �������S� C�_�g�y��������� ӏ�����7�a��� ���ﲟ���ӟ� ��0��T�?�x�c�u� ����ү������,� #�P��_t�������	� ���o���(��L� ^�pς�AϦϸ����� �� ��$���H�Z�l� ~�=ߢߴ����ߗ��� � ���D�V�h�z�9� ����������
�� ��@�R�d�v�5����� ����������< N`r1����? ��8J\ n-������ �/�4/F/X/j/)/ �/�/�/�/�/�/�/? oc�9?Q�]?M?i?q? �?�?�?�?�?�?OO O%O7OkO[OwOO�O �O�O�O�O�O�O_C_ 3_O_W_i_�_�_�_�_ �_�_�_oo'oQoAo uou�?�o�o�o�o�o �o D/Aze �������� �@�7�d�v��/���� ��Џ/�􏃏�*�<� N��r�����U���̟ ޟ🯟�&�8�J�	� n�����Q���ȯگ� ���"�4�F��j�|� ��M���Ŀֿ迧�� �0�B��f�xϊ�I� �������ϣ���,� >���b�t߆�Eߖ߼� �������(�:�� ^�p��A������� �� ��$�6���Z�l� ~�=�������������  2)?MeoYa s������ '[Kgo� �������3/ #/?/G/Y/�/}/�/�/ �/�/�/�/�/?A?1?�e?U?q?y?�1�$P�LCL_GRP �1���1�� D�0��?�  �6s��?~5?�:�0� O�:O%O^OIO�OmO O�O�O�O�O _�O�= 1_�OX_�O|_g_�_�_ �_�_�_�_�_o	oBo )o#_uo7o�o3o�o�o �o�o�o>)b M�mgo�{�w ��(��8�^�I����m�����ʏ<	�$VCAX_REF�0� 2�5� t 
 ����EREN/CE 1��׏7��I�[�m�������2 �ԟ���
��.�@����3ß|������� į֯�S��4k�$� 6�H�Z�l�~������5�̿޿���&� 8ϣ���4��zόϞ� �������ϱ�7c�� .�@�R�d�v߈����8�����������0���9��l�~���������C�FA�CTORY DATA\��'�9�K�]�o������9�������������	 `��GYk
�2_� ��������2_�Pbt ����'j�?� 
//./@/R/d/'� ��/�/�/�/�/�/? '���/H?Z?l?~?�? �?�?'b�7?�?OO &O8OJO\O'
��?�O �O�O�O�O�O_'�� �O@_R_d_v_�_�_�_ 'Z�/_�_�_oo0o BoTo���_�o�o�o�o �o�o�o��/A Sew%�����3��%�7�I�[� m���_�t7��Ώ�� ���(������d� v���������П;��� �/��0�B�T�f�x� 㟥�/?��Ưد��� � ������?\�n��� ������ȿ3���O� �(�:�L�^�p�ۿ�� '_�Ͼ��������� �ϥ��_T�f�xߊߜ� ����_oqo����,� >�P�b�t����� ��������(�:�L����4��������� ������*�p���0B Tfx��S� ��� 2D� �������� �W��(/:/L/^/ p/�/�/�K��/�/ �/??*?<?�/� x?�?�?�?�?�?�?O? �� O2ODOVOhOzO �O�?C��O�O�O�O _"_4_����j_|_�_ �_�_�_�_�_��	�o !o3oEoWoio��o�o �o�d